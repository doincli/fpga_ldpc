module error_comp(
    clk    ,
    rst_n  ,
    r_en  ,
    data_in,
    H_in,
    data_out
    );

    //��������
    parameter      DATA_W =         256;
    parameter      DATA_H_in =         4096;

    //�����źŶ���
    input               clk    ;
    input               rst_n  ;
    input[DATA_W-1:0]  data_in ;
    input[DATA_H_in-1:0]   H_in   ;
    input    r_en              ;

    //����źŶ���
    output [15:0]  data_out;

    //����ź�reg����
    reg   [15:0]  data_out   ;

    wire add_cnt;
    wire end_cnt;
    reg [1:0] cnt;
    always @(posedge clk or negedge rst_n)begin
        if(!rst_n)begin
            cnt <= 0;
        end
        else if(add_cnt)begin
            if(end_cnt)
                cnt <= 0;
            else
                cnt <= cnt + 1;
        end
    end

    assign add_cnt = r_en==1;       
    assign end_cnt = add_cnt && cnt==1 ;   

     //����ͼ���ļ���
     always  @(posedge clk or negedge rst_n)begin
         if(rst_n==1'b0)begin
               data_out <= 0 ;
         end
         else if(r_en==0&&cnt==0)begin
         data_out[0]<=(data_in[0]&H_in[0])^(data_in[1]&H_in[1])^(data_in[2]&H_in[2])^(data_in[3]&H_in[3])^(data_in[4]&H_in[4])^(data_in[5]&H_in[5])^(data_in[6]&H_in[6])^(data_in[7]&H_in[7])^(data_in[8]&H_in[8])^(data_in[9]&H_in[9])^(data_in[10]&H_in[10])^(data_in[11]&H_in[11])^(data_in[12]&H_in[12])^(data_in[13]&H_in[13])^(data_in[14]&H_in[14])^(data_in[15]&H_in[15])^(data_in[16]&H_in[16])^(data_in[17]&H_in[17])^(data_in[18]&H_in[18])^(data_in[19]&H_in[19])^(data_in[20]&H_in[20])^(data_in[21]&H_in[21])^(data_in[22]&H_in[22])^(data_in[23]&H_in[23])^(data_in[24]&H_in[24])^(data_in[25]&H_in[25])^(data_in[26]&H_in[26])^(data_in[27]&H_in[27])^(data_in[28]&H_in[28])^(data_in[29]&H_in[29])^(data_in[30]&H_in[30])^(data_in[31]&H_in[31])^(data_in[32]&H_in[32])^(data_in[33]&H_in[33])^(data_in[34]&H_in[34])^(data_in[35]&H_in[35])^(data_in[36]&H_in[36])^(data_in[37]&H_in[37])^(data_in[38]&H_in[38])^(data_in[39]&H_in[39])^(data_in[40]&H_in[40])^(data_in[41]&H_in[41])^(data_in[42]&H_in[42])^(data_in[43]&H_in[43])^(data_in[44]&H_in[44])^(data_in[45]&H_in[45])^(data_in[46]&H_in[46])^(data_in[47]&H_in[47])^(data_in[48]&H_in[48])^(data_in[49]&H_in[49])^(data_in[50]&H_in[50])^(data_in[51]&H_in[51])^(data_in[52]&H_in[52])^(data_in[53]&H_in[53])^(data_in[54]&H_in[54])^(data_in[55]&H_in[55])^(data_in[56]&H_in[56])^(data_in[57]&H_in[57])^(data_in[58]&H_in[58])^(data_in[59]&H_in[59])^(data_in[60]&H_in[60])^(data_in[61]&H_in[61])^(data_in[62]&H_in[62])^(data_in[63]&H_in[63])^(data_in[64]&H_in[64])^(data_in[65]&H_in[65])^(data_in[66]&H_in[66])^(data_in[67]&H_in[67])^(data_in[68]&H_in[68])^(data_in[69]&H_in[69])^(data_in[70]&H_in[70])^(data_in[71]&H_in[71])^(data_in[72]&H_in[72])^(data_in[73]&H_in[73])^(data_in[74]&H_in[74])^(data_in[75]&H_in[75])^(data_in[76]&H_in[76])^(data_in[77]&H_in[77])^(data_in[78]&H_in[78])^(data_in[79]&H_in[79])^(data_in[80]&H_in[80])^(data_in[81]&H_in[81])^(data_in[82]&H_in[82])^(data_in[83]&H_in[83])^(data_in[84]&H_in[84])^(data_in[85]&H_in[85])^(data_in[86]&H_in[86])^(data_in[87]&H_in[87])^(data_in[88]&H_in[88])^(data_in[89]&H_in[89])^(data_in[90]&H_in[90])^(data_in[91]&H_in[91])^(data_in[92]&H_in[92])^(data_in[93]&H_in[93])^(data_in[94]&H_in[94])^(data_in[95]&H_in[95])^(data_in[96]&H_in[96])^(data_in[97]&H_in[97])^(data_in[98]&H_in[98])^(data_in[99]&H_in[99])^(data_in[100]&H_in[100])^(data_in[101]&H_in[101])^(data_in[102]&H_in[102])^(data_in[103]&H_in[103])^(data_in[104]&H_in[104])^(data_in[105]&H_in[105])^(data_in[106]&H_in[106])^(data_in[107]&H_in[107])^(data_in[108]&H_in[108])^(data_in[109]&H_in[109])^(data_in[110]&H_in[110])^(data_in[111]&H_in[111])^(data_in[112]&H_in[112])^(data_in[113]&H_in[113])^(data_in[114]&H_in[114])^(data_in[115]&H_in[115])^(data_in[116]&H_in[116])^(data_in[117]&H_in[117])^(data_in[118]&H_in[118])^(data_in[119]&H_in[119])^(data_in[120]&H_in[120])^(data_in[121]&H_in[121])^(data_in[122]&H_in[122])^(data_in[123]&H_in[123])^(data_in[124]&H_in[124])^(data_in[125]&H_in[125])^(data_in[126]&H_in[126])^(data_in[127]&H_in[127])^(data_in[128]&H_in[128])^(data_in[129]&H_in[129])^(data_in[130]&H_in[130])^(data_in[131]&H_in[131])^(data_in[132]&H_in[132])^(data_in[133]&H_in[133])^(data_in[134]&H_in[134])^(data_in[135]&H_in[135])^(data_in[136]&H_in[136])^(data_in[137]&H_in[137])^(data_in[138]&H_in[138])^(data_in[139]&H_in[139])^(data_in[140]&H_in[140])^(data_in[141]&H_in[141])^(data_in[142]&H_in[142])^(data_in[143]&H_in[143])^(data_in[144]&H_in[144])^(data_in[145]&H_in[145])^(data_in[146]&H_in[146])^(data_in[147]&H_in[147])^(data_in[148]&H_in[148])^(data_in[149]&H_in[149])^(data_in[150]&H_in[150])^(data_in[151]&H_in[151])^(data_in[152]&H_in[152])^(data_in[153]&H_in[153])^(data_in[154]&H_in[154])^(data_in[155]&H_in[155])^(data_in[156]&H_in[156])^(data_in[157]&H_in[157])^(data_in[158]&H_in[158])^(data_in[159]&H_in[159])^(data_in[160]&H_in[160])^(data_in[161]&H_in[161])^(data_in[162]&H_in[162])^(data_in[163]&H_in[163])^(data_in[164]&H_in[164])^(data_in[165]&H_in[165])^(data_in[166]&H_in[166])^(data_in[167]&H_in[167])^(data_in[168]&H_in[168])^(data_in[169]&H_in[169])^(data_in[170]&H_in[170])^(data_in[171]&H_in[171])^(data_in[172]&H_in[172])^(data_in[173]&H_in[173])^(data_in[174]&H_in[174])^(data_in[175]&H_in[175])^(data_in[176]&H_in[176])^(data_in[177]&H_in[177])^(data_in[178]&H_in[178])^(data_in[179]&H_in[179])^(data_in[180]&H_in[180])^(data_in[181]&H_in[181])^(data_in[182]&H_in[182])^(data_in[183]&H_in[183])^(data_in[184]&H_in[184])^(data_in[185]&H_in[185])^(data_in[186]&H_in[186])^(data_in[187]&H_in[187])^(data_in[188]&H_in[188])^(data_in[189]&H_in[189])^(data_in[190]&H_in[190])^(data_in[191]&H_in[191])^(data_in[192]&H_in[192])^(data_in[193]&H_in[193])^(data_in[194]&H_in[194])^(data_in[195]&H_in[195])^(data_in[196]&H_in[196])^(data_in[197]&H_in[197])^(data_in[198]&H_in[198])^(data_in[199]&H_in[199])^(data_in[200]&H_in[200])^(data_in[201]&H_in[201])^(data_in[202]&H_in[202])^(data_in[203]&H_in[203])^(data_in[204]&H_in[204])^(data_in[205]&H_in[205])^(data_in[206]&H_in[206])^(data_in[207]&H_in[207])^(data_in[208]&H_in[208])^(data_in[209]&H_in[209])^(data_in[210]&H_in[210])^(data_in[211]&H_in[211])^(data_in[212]&H_in[212])^(data_in[213]&H_in[213])^(data_in[214]&H_in[214])^(data_in[215]&H_in[215])^(data_in[216]&H_in[216])^(data_in[217]&H_in[217])^(data_in[218]&H_in[218])^(data_in[219]&H_in[219])^(data_in[220]&H_in[220])^(data_in[221]&H_in[221])^(data_in[222]&H_in[222])^(data_in[223]&H_in[223])^(data_in[224]&H_in[224])^(data_in[225]&H_in[225])^(data_in[226]&H_in[226])^(data_in[227]&H_in[227])^(data_in[228]&H_in[228])^(data_in[229]&H_in[229])^(data_in[230]&H_in[230])^(data_in[231]&H_in[231])^(data_in[232]&H_in[232])^(data_in[233]&H_in[233])^(data_in[234]&H_in[234])^(data_in[235]&H_in[235])^(data_in[236]&H_in[236])^(data_in[237]&H_in[237])^(data_in[238]&H_in[238])^(data_in[239]&H_in[239])^(data_in[240]&H_in[240])^(data_in[241]&H_in[241])^(data_in[242]&H_in[242])^(data_in[243]&H_in[243])^(data_in[244]&H_in[244])^(data_in[245]&H_in[245])^(data_in[246]&H_in[246])^(data_in[247]&H_in[247])^(data_in[248]&H_in[248])^(data_in[249]&H_in[249])^(data_in[250]&H_in[250])^(data_in[251]&H_in[251])^(data_in[252]&H_in[252])^(data_in[253]&H_in[253])^(data_in[254]&H_in[254])^(data_in[255]&H_in[255]);
         data_out[1]<=(data_in[0]&H_in[256])^(data_in[1]&H_in[257])^(data_in[2]&H_in[258])^(data_in[3]&H_in[259])^(data_in[4]&H_in[260])^(data_in[5]&H_in[261])^(data_in[6]&H_in[262])^(data_in[7]&H_in[263])^(data_in[8]&H_in[264])^(data_in[9]&H_in[265])^(data_in[10]&H_in[266])^(data_in[11]&H_in[267])^(data_in[12]&H_in[268])^(data_in[13]&H_in[269])^(data_in[14]&H_in[270])^(data_in[15]&H_in[271])^(data_in[16]&H_in[272])^(data_in[17]&H_in[273])^(data_in[18]&H_in[274])^(data_in[19]&H_in[275])^(data_in[20]&H_in[276])^(data_in[21]&H_in[277])^(data_in[22]&H_in[278])^(data_in[23]&H_in[279])^(data_in[24]&H_in[280])^(data_in[25]&H_in[281])^(data_in[26]&H_in[282])^(data_in[27]&H_in[283])^(data_in[28]&H_in[284])^(data_in[29]&H_in[285])^(data_in[30]&H_in[286])^(data_in[31]&H_in[287])^(data_in[32]&H_in[288])^(data_in[33]&H_in[289])^(data_in[34]&H_in[290])^(data_in[35]&H_in[291])^(data_in[36]&H_in[292])^(data_in[37]&H_in[293])^(data_in[38]&H_in[294])^(data_in[39]&H_in[295])^(data_in[40]&H_in[296])^(data_in[41]&H_in[297])^(data_in[42]&H_in[298])^(data_in[43]&H_in[299])^(data_in[44]&H_in[300])^(data_in[45]&H_in[301])^(data_in[46]&H_in[302])^(data_in[47]&H_in[303])^(data_in[48]&H_in[304])^(data_in[49]&H_in[305])^(data_in[50]&H_in[306])^(data_in[51]&H_in[307])^(data_in[52]&H_in[308])^(data_in[53]&H_in[309])^(data_in[54]&H_in[310])^(data_in[55]&H_in[311])^(data_in[56]&H_in[312])^(data_in[57]&H_in[313])^(data_in[58]&H_in[314])^(data_in[59]&H_in[315])^(data_in[60]&H_in[316])^(data_in[61]&H_in[317])^(data_in[62]&H_in[318])^(data_in[63]&H_in[319])^(data_in[64]&H_in[320])^(data_in[65]&H_in[321])^(data_in[66]&H_in[322])^(data_in[67]&H_in[323])^(data_in[68]&H_in[324])^(data_in[69]&H_in[325])^(data_in[70]&H_in[326])^(data_in[71]&H_in[327])^(data_in[72]&H_in[328])^(data_in[73]&H_in[329])^(data_in[74]&H_in[330])^(data_in[75]&H_in[331])^(data_in[76]&H_in[332])^(data_in[77]&H_in[333])^(data_in[78]&H_in[334])^(data_in[79]&H_in[335])^(data_in[80]&H_in[336])^(data_in[81]&H_in[337])^(data_in[82]&H_in[338])^(data_in[83]&H_in[339])^(data_in[84]&H_in[340])^(data_in[85]&H_in[341])^(data_in[86]&H_in[342])^(data_in[87]&H_in[343])^(data_in[88]&H_in[344])^(data_in[89]&H_in[345])^(data_in[90]&H_in[346])^(data_in[91]&H_in[347])^(data_in[92]&H_in[348])^(data_in[93]&H_in[349])^(data_in[94]&H_in[350])^(data_in[95]&H_in[351])^(data_in[96]&H_in[352])^(data_in[97]&H_in[353])^(data_in[98]&H_in[354])^(data_in[99]&H_in[355])^(data_in[100]&H_in[356])^(data_in[101]&H_in[357])^(data_in[102]&H_in[358])^(data_in[103]&H_in[359])^(data_in[104]&H_in[360])^(data_in[105]&H_in[361])^(data_in[106]&H_in[362])^(data_in[107]&H_in[363])^(data_in[108]&H_in[364])^(data_in[109]&H_in[365])^(data_in[110]&H_in[366])^(data_in[111]&H_in[367])^(data_in[112]&H_in[368])^(data_in[113]&H_in[369])^(data_in[114]&H_in[370])^(data_in[115]&H_in[371])^(data_in[116]&H_in[372])^(data_in[117]&H_in[373])^(data_in[118]&H_in[374])^(data_in[119]&H_in[375])^(data_in[120]&H_in[376])^(data_in[121]&H_in[377])^(data_in[122]&H_in[378])^(data_in[123]&H_in[379])^(data_in[124]&H_in[380])^(data_in[125]&H_in[381])^(data_in[126]&H_in[382])^(data_in[127]&H_in[383])^(data_in[128]&H_in[384])^(data_in[129]&H_in[385])^(data_in[130]&H_in[386])^(data_in[131]&H_in[387])^(data_in[132]&H_in[388])^(data_in[133]&H_in[389])^(data_in[134]&H_in[390])^(data_in[135]&H_in[391])^(data_in[136]&H_in[392])^(data_in[137]&H_in[393])^(data_in[138]&H_in[394])^(data_in[139]&H_in[395])^(data_in[140]&H_in[396])^(data_in[141]&H_in[397])^(data_in[142]&H_in[398])^(data_in[143]&H_in[399])^(data_in[144]&H_in[400])^(data_in[145]&H_in[401])^(data_in[146]&H_in[402])^(data_in[147]&H_in[403])^(data_in[148]&H_in[404])^(data_in[149]&H_in[405])^(data_in[150]&H_in[406])^(data_in[151]&H_in[407])^(data_in[152]&H_in[408])^(data_in[153]&H_in[409])^(data_in[154]&H_in[410])^(data_in[155]&H_in[411])^(data_in[156]&H_in[412])^(data_in[157]&H_in[413])^(data_in[158]&H_in[414])^(data_in[159]&H_in[415])^(data_in[160]&H_in[416])^(data_in[161]&H_in[417])^(data_in[162]&H_in[418])^(data_in[163]&H_in[419])^(data_in[164]&H_in[420])^(data_in[165]&H_in[421])^(data_in[166]&H_in[422])^(data_in[167]&H_in[423])^(data_in[168]&H_in[424])^(data_in[169]&H_in[425])^(data_in[170]&H_in[426])^(data_in[171]&H_in[427])^(data_in[172]&H_in[428])^(data_in[173]&H_in[429])^(data_in[174]&H_in[430])^(data_in[175]&H_in[431])^(data_in[176]&H_in[432])^(data_in[177]&H_in[433])^(data_in[178]&H_in[434])^(data_in[179]&H_in[435])^(data_in[180]&H_in[436])^(data_in[181]&H_in[437])^(data_in[182]&H_in[438])^(data_in[183]&H_in[439])^(data_in[184]&H_in[440])^(data_in[185]&H_in[441])^(data_in[186]&H_in[442])^(data_in[187]&H_in[443])^(data_in[188]&H_in[444])^(data_in[189]&H_in[445])^(data_in[190]&H_in[446])^(data_in[191]&H_in[447])^(data_in[192]&H_in[448])^(data_in[193]&H_in[449])^(data_in[194]&H_in[450])^(data_in[195]&H_in[451])^(data_in[196]&H_in[452])^(data_in[197]&H_in[453])^(data_in[198]&H_in[454])^(data_in[199]&H_in[455])^(data_in[200]&H_in[456])^(data_in[201]&H_in[457])^(data_in[202]&H_in[458])^(data_in[203]&H_in[459])^(data_in[204]&H_in[460])^(data_in[205]&H_in[461])^(data_in[206]&H_in[462])^(data_in[207]&H_in[463])^(data_in[208]&H_in[464])^(data_in[209]&H_in[465])^(data_in[210]&H_in[466])^(data_in[211]&H_in[467])^(data_in[212]&H_in[468])^(data_in[213]&H_in[469])^(data_in[214]&H_in[470])^(data_in[215]&H_in[471])^(data_in[216]&H_in[472])^(data_in[217]&H_in[473])^(data_in[218]&H_in[474])^(data_in[219]&H_in[475])^(data_in[220]&H_in[476])^(data_in[221]&H_in[477])^(data_in[222]&H_in[478])^(data_in[223]&H_in[479])^(data_in[224]&H_in[480])^(data_in[225]&H_in[481])^(data_in[226]&H_in[482])^(data_in[227]&H_in[483])^(data_in[228]&H_in[484])^(data_in[229]&H_in[485])^(data_in[230]&H_in[486])^(data_in[231]&H_in[487])^(data_in[232]&H_in[488])^(data_in[233]&H_in[489])^(data_in[234]&H_in[490])^(data_in[235]&H_in[491])^(data_in[236]&H_in[492])^(data_in[237]&H_in[493])^(data_in[238]&H_in[494])^(data_in[239]&H_in[495])^(data_in[240]&H_in[496])^(data_in[241]&H_in[497])^(data_in[242]&H_in[498])^(data_in[243]&H_in[499])^(data_in[244]&H_in[500])^(data_in[245]&H_in[501])^(data_in[246]&H_in[502])^(data_in[247]&H_in[503])^(data_in[248]&H_in[504])^(data_in[249]&H_in[505])^(data_in[250]&H_in[506])^(data_in[251]&H_in[507])^(data_in[252]&H_in[508])^(data_in[253]&H_in[509])^(data_in[254]&H_in[510])^(data_in[255]&H_in[511]);
         data_out[2]<=(data_in[0]&H_in[512])^(data_in[1]&H_in[513])^(data_in[2]&H_in[514])^(data_in[3]&H_in[515])^(data_in[4]&H_in[516])^(data_in[5]&H_in[517])^(data_in[6]&H_in[518])^(data_in[7]&H_in[519])^(data_in[8]&H_in[520])^(data_in[9]&H_in[521])^(data_in[10]&H_in[522])^(data_in[11]&H_in[523])^(data_in[12]&H_in[524])^(data_in[13]&H_in[525])^(data_in[14]&H_in[526])^(data_in[15]&H_in[527])^(data_in[16]&H_in[528])^(data_in[17]&H_in[529])^(data_in[18]&H_in[530])^(data_in[19]&H_in[531])^(data_in[20]&H_in[532])^(data_in[21]&H_in[533])^(data_in[22]&H_in[534])^(data_in[23]&H_in[535])^(data_in[24]&H_in[536])^(data_in[25]&H_in[537])^(data_in[26]&H_in[538])^(data_in[27]&H_in[539])^(data_in[28]&H_in[540])^(data_in[29]&H_in[541])^(data_in[30]&H_in[542])^(data_in[31]&H_in[543])^(data_in[32]&H_in[544])^(data_in[33]&H_in[545])^(data_in[34]&H_in[546])^(data_in[35]&H_in[547])^(data_in[36]&H_in[548])^(data_in[37]&H_in[549])^(data_in[38]&H_in[550])^(data_in[39]&H_in[551])^(data_in[40]&H_in[552])^(data_in[41]&H_in[553])^(data_in[42]&H_in[554])^(data_in[43]&H_in[555])^(data_in[44]&H_in[556])^(data_in[45]&H_in[557])^(data_in[46]&H_in[558])^(data_in[47]&H_in[559])^(data_in[48]&H_in[560])^(data_in[49]&H_in[561])^(data_in[50]&H_in[562])^(data_in[51]&H_in[563])^(data_in[52]&H_in[564])^(data_in[53]&H_in[565])^(data_in[54]&H_in[566])^(data_in[55]&H_in[567])^(data_in[56]&H_in[568])^(data_in[57]&H_in[569])^(data_in[58]&H_in[570])^(data_in[59]&H_in[571])^(data_in[60]&H_in[572])^(data_in[61]&H_in[573])^(data_in[62]&H_in[574])^(data_in[63]&H_in[575])^(data_in[64]&H_in[576])^(data_in[65]&H_in[577])^(data_in[66]&H_in[578])^(data_in[67]&H_in[579])^(data_in[68]&H_in[580])^(data_in[69]&H_in[581])^(data_in[70]&H_in[582])^(data_in[71]&H_in[583])^(data_in[72]&H_in[584])^(data_in[73]&H_in[585])^(data_in[74]&H_in[586])^(data_in[75]&H_in[587])^(data_in[76]&H_in[588])^(data_in[77]&H_in[589])^(data_in[78]&H_in[590])^(data_in[79]&H_in[591])^(data_in[80]&H_in[592])^(data_in[81]&H_in[593])^(data_in[82]&H_in[594])^(data_in[83]&H_in[595])^(data_in[84]&H_in[596])^(data_in[85]&H_in[597])^(data_in[86]&H_in[598])^(data_in[87]&H_in[599])^(data_in[88]&H_in[600])^(data_in[89]&H_in[601])^(data_in[90]&H_in[602])^(data_in[91]&H_in[603])^(data_in[92]&H_in[604])^(data_in[93]&H_in[605])^(data_in[94]&H_in[606])^(data_in[95]&H_in[607])^(data_in[96]&H_in[608])^(data_in[97]&H_in[609])^(data_in[98]&H_in[610])^(data_in[99]&H_in[611])^(data_in[100]&H_in[612])^(data_in[101]&H_in[613])^(data_in[102]&H_in[614])^(data_in[103]&H_in[615])^(data_in[104]&H_in[616])^(data_in[105]&H_in[617])^(data_in[106]&H_in[618])^(data_in[107]&H_in[619])^(data_in[108]&H_in[620])^(data_in[109]&H_in[621])^(data_in[110]&H_in[622])^(data_in[111]&H_in[623])^(data_in[112]&H_in[624])^(data_in[113]&H_in[625])^(data_in[114]&H_in[626])^(data_in[115]&H_in[627])^(data_in[116]&H_in[628])^(data_in[117]&H_in[629])^(data_in[118]&H_in[630])^(data_in[119]&H_in[631])^(data_in[120]&H_in[632])^(data_in[121]&H_in[633])^(data_in[122]&H_in[634])^(data_in[123]&H_in[635])^(data_in[124]&H_in[636])^(data_in[125]&H_in[637])^(data_in[126]&H_in[638])^(data_in[127]&H_in[639])^(data_in[128]&H_in[640])^(data_in[129]&H_in[641])^(data_in[130]&H_in[642])^(data_in[131]&H_in[643])^(data_in[132]&H_in[644])^(data_in[133]&H_in[645])^(data_in[134]&H_in[646])^(data_in[135]&H_in[647])^(data_in[136]&H_in[648])^(data_in[137]&H_in[649])^(data_in[138]&H_in[650])^(data_in[139]&H_in[651])^(data_in[140]&H_in[652])^(data_in[141]&H_in[653])^(data_in[142]&H_in[654])^(data_in[143]&H_in[655])^(data_in[144]&H_in[656])^(data_in[145]&H_in[657])^(data_in[146]&H_in[658])^(data_in[147]&H_in[659])^(data_in[148]&H_in[660])^(data_in[149]&H_in[661])^(data_in[150]&H_in[662])^(data_in[151]&H_in[663])^(data_in[152]&H_in[664])^(data_in[153]&H_in[665])^(data_in[154]&H_in[666])^(data_in[155]&H_in[667])^(data_in[156]&H_in[668])^(data_in[157]&H_in[669])^(data_in[158]&H_in[670])^(data_in[159]&H_in[671])^(data_in[160]&H_in[672])^(data_in[161]&H_in[673])^(data_in[162]&H_in[674])^(data_in[163]&H_in[675])^(data_in[164]&H_in[676])^(data_in[165]&H_in[677])^(data_in[166]&H_in[678])^(data_in[167]&H_in[679])^(data_in[168]&H_in[680])^(data_in[169]&H_in[681])^(data_in[170]&H_in[682])^(data_in[171]&H_in[683])^(data_in[172]&H_in[684])^(data_in[173]&H_in[685])^(data_in[174]&H_in[686])^(data_in[175]&H_in[687])^(data_in[176]&H_in[688])^(data_in[177]&H_in[689])^(data_in[178]&H_in[690])^(data_in[179]&H_in[691])^(data_in[180]&H_in[692])^(data_in[181]&H_in[693])^(data_in[182]&H_in[694])^(data_in[183]&H_in[695])^(data_in[184]&H_in[696])^(data_in[185]&H_in[697])^(data_in[186]&H_in[698])^(data_in[187]&H_in[699])^(data_in[188]&H_in[700])^(data_in[189]&H_in[701])^(data_in[190]&H_in[702])^(data_in[191]&H_in[703])^(data_in[192]&H_in[704])^(data_in[193]&H_in[705])^(data_in[194]&H_in[706])^(data_in[195]&H_in[707])^(data_in[196]&H_in[708])^(data_in[197]&H_in[709])^(data_in[198]&H_in[710])^(data_in[199]&H_in[711])^(data_in[200]&H_in[712])^(data_in[201]&H_in[713])^(data_in[202]&H_in[714])^(data_in[203]&H_in[715])^(data_in[204]&H_in[716])^(data_in[205]&H_in[717])^(data_in[206]&H_in[718])^(data_in[207]&H_in[719])^(data_in[208]&H_in[720])^(data_in[209]&H_in[721])^(data_in[210]&H_in[722])^(data_in[211]&H_in[723])^(data_in[212]&H_in[724])^(data_in[213]&H_in[725])^(data_in[214]&H_in[726])^(data_in[215]&H_in[727])^(data_in[216]&H_in[728])^(data_in[217]&H_in[729])^(data_in[218]&H_in[730])^(data_in[219]&H_in[731])^(data_in[220]&H_in[732])^(data_in[221]&H_in[733])^(data_in[222]&H_in[734])^(data_in[223]&H_in[735])^(data_in[224]&H_in[736])^(data_in[225]&H_in[737])^(data_in[226]&H_in[738])^(data_in[227]&H_in[739])^(data_in[228]&H_in[740])^(data_in[229]&H_in[741])^(data_in[230]&H_in[742])^(data_in[231]&H_in[743])^(data_in[232]&H_in[744])^(data_in[233]&H_in[745])^(data_in[234]&H_in[746])^(data_in[235]&H_in[747])^(data_in[236]&H_in[748])^(data_in[237]&H_in[749])^(data_in[238]&H_in[750])^(data_in[239]&H_in[751])^(data_in[240]&H_in[752])^(data_in[241]&H_in[753])^(data_in[242]&H_in[754])^(data_in[243]&H_in[755])^(data_in[244]&H_in[756])^(data_in[245]&H_in[757])^(data_in[246]&H_in[758])^(data_in[247]&H_in[759])^(data_in[248]&H_in[760])^(data_in[249]&H_in[761])^(data_in[250]&H_in[762])^(data_in[251]&H_in[763])^(data_in[252]&H_in[764])^(data_in[253]&H_in[765])^(data_in[254]&H_in[766])^(data_in[255]&H_in[767]);
         data_out[3]<=(data_in[0]&H_in[768])^(data_in[1]&H_in[769])^(data_in[2]&H_in[770])^(data_in[3]&H_in[771])^(data_in[4]&H_in[772])^(data_in[5]&H_in[773])^(data_in[6]&H_in[774])^(data_in[7]&H_in[775])^(data_in[8]&H_in[776])^(data_in[9]&H_in[777])^(data_in[10]&H_in[778])^(data_in[11]&H_in[779])^(data_in[12]&H_in[780])^(data_in[13]&H_in[781])^(data_in[14]&H_in[782])^(data_in[15]&H_in[783])^(data_in[16]&H_in[784])^(data_in[17]&H_in[785])^(data_in[18]&H_in[786])^(data_in[19]&H_in[787])^(data_in[20]&H_in[788])^(data_in[21]&H_in[789])^(data_in[22]&H_in[790])^(data_in[23]&H_in[791])^(data_in[24]&H_in[792])^(data_in[25]&H_in[793])^(data_in[26]&H_in[794])^(data_in[27]&H_in[795])^(data_in[28]&H_in[796])^(data_in[29]&H_in[797])^(data_in[30]&H_in[798])^(data_in[31]&H_in[799])^(data_in[32]&H_in[800])^(data_in[33]&H_in[801])^(data_in[34]&H_in[802])^(data_in[35]&H_in[803])^(data_in[36]&H_in[804])^(data_in[37]&H_in[805])^(data_in[38]&H_in[806])^(data_in[39]&H_in[807])^(data_in[40]&H_in[808])^(data_in[41]&H_in[809])^(data_in[42]&H_in[810])^(data_in[43]&H_in[811])^(data_in[44]&H_in[812])^(data_in[45]&H_in[813])^(data_in[46]&H_in[814])^(data_in[47]&H_in[815])^(data_in[48]&H_in[816])^(data_in[49]&H_in[817])^(data_in[50]&H_in[818])^(data_in[51]&H_in[819])^(data_in[52]&H_in[820])^(data_in[53]&H_in[821])^(data_in[54]&H_in[822])^(data_in[55]&H_in[823])^(data_in[56]&H_in[824])^(data_in[57]&H_in[825])^(data_in[58]&H_in[826])^(data_in[59]&H_in[827])^(data_in[60]&H_in[828])^(data_in[61]&H_in[829])^(data_in[62]&H_in[830])^(data_in[63]&H_in[831])^(data_in[64]&H_in[832])^(data_in[65]&H_in[833])^(data_in[66]&H_in[834])^(data_in[67]&H_in[835])^(data_in[68]&H_in[836])^(data_in[69]&H_in[837])^(data_in[70]&H_in[838])^(data_in[71]&H_in[839])^(data_in[72]&H_in[840])^(data_in[73]&H_in[841])^(data_in[74]&H_in[842])^(data_in[75]&H_in[843])^(data_in[76]&H_in[844])^(data_in[77]&H_in[845])^(data_in[78]&H_in[846])^(data_in[79]&H_in[847])^(data_in[80]&H_in[848])^(data_in[81]&H_in[849])^(data_in[82]&H_in[850])^(data_in[83]&H_in[851])^(data_in[84]&H_in[852])^(data_in[85]&H_in[853])^(data_in[86]&H_in[854])^(data_in[87]&H_in[855])^(data_in[88]&H_in[856])^(data_in[89]&H_in[857])^(data_in[90]&H_in[858])^(data_in[91]&H_in[859])^(data_in[92]&H_in[860])^(data_in[93]&H_in[861])^(data_in[94]&H_in[862])^(data_in[95]&H_in[863])^(data_in[96]&H_in[864])^(data_in[97]&H_in[865])^(data_in[98]&H_in[866])^(data_in[99]&H_in[867])^(data_in[100]&H_in[868])^(data_in[101]&H_in[869])^(data_in[102]&H_in[870])^(data_in[103]&H_in[871])^(data_in[104]&H_in[872])^(data_in[105]&H_in[873])^(data_in[106]&H_in[874])^(data_in[107]&H_in[875])^(data_in[108]&H_in[876])^(data_in[109]&H_in[877])^(data_in[110]&H_in[878])^(data_in[111]&H_in[879])^(data_in[112]&H_in[880])^(data_in[113]&H_in[881])^(data_in[114]&H_in[882])^(data_in[115]&H_in[883])^(data_in[116]&H_in[884])^(data_in[117]&H_in[885])^(data_in[118]&H_in[886])^(data_in[119]&H_in[887])^(data_in[120]&H_in[888])^(data_in[121]&H_in[889])^(data_in[122]&H_in[890])^(data_in[123]&H_in[891])^(data_in[124]&H_in[892])^(data_in[125]&H_in[893])^(data_in[126]&H_in[894])^(data_in[127]&H_in[895])^(data_in[128]&H_in[896])^(data_in[129]&H_in[897])^(data_in[130]&H_in[898])^(data_in[131]&H_in[899])^(data_in[132]&H_in[900])^(data_in[133]&H_in[901])^(data_in[134]&H_in[902])^(data_in[135]&H_in[903])^(data_in[136]&H_in[904])^(data_in[137]&H_in[905])^(data_in[138]&H_in[906])^(data_in[139]&H_in[907])^(data_in[140]&H_in[908])^(data_in[141]&H_in[909])^(data_in[142]&H_in[910])^(data_in[143]&H_in[911])^(data_in[144]&H_in[912])^(data_in[145]&H_in[913])^(data_in[146]&H_in[914])^(data_in[147]&H_in[915])^(data_in[148]&H_in[916])^(data_in[149]&H_in[917])^(data_in[150]&H_in[918])^(data_in[151]&H_in[919])^(data_in[152]&H_in[920])^(data_in[153]&H_in[921])^(data_in[154]&H_in[922])^(data_in[155]&H_in[923])^(data_in[156]&H_in[924])^(data_in[157]&H_in[925])^(data_in[158]&H_in[926])^(data_in[159]&H_in[927])^(data_in[160]&H_in[928])^(data_in[161]&H_in[929])^(data_in[162]&H_in[930])^(data_in[163]&H_in[931])^(data_in[164]&H_in[932])^(data_in[165]&H_in[933])^(data_in[166]&H_in[934])^(data_in[167]&H_in[935])^(data_in[168]&H_in[936])^(data_in[169]&H_in[937])^(data_in[170]&H_in[938])^(data_in[171]&H_in[939])^(data_in[172]&H_in[940])^(data_in[173]&H_in[941])^(data_in[174]&H_in[942])^(data_in[175]&H_in[943])^(data_in[176]&H_in[944])^(data_in[177]&H_in[945])^(data_in[178]&H_in[946])^(data_in[179]&H_in[947])^(data_in[180]&H_in[948])^(data_in[181]&H_in[949])^(data_in[182]&H_in[950])^(data_in[183]&H_in[951])^(data_in[184]&H_in[952])^(data_in[185]&H_in[953])^(data_in[186]&H_in[954])^(data_in[187]&H_in[955])^(data_in[188]&H_in[956])^(data_in[189]&H_in[957])^(data_in[190]&H_in[958])^(data_in[191]&H_in[959])^(data_in[192]&H_in[960])^(data_in[193]&H_in[961])^(data_in[194]&H_in[962])^(data_in[195]&H_in[963])^(data_in[196]&H_in[964])^(data_in[197]&H_in[965])^(data_in[198]&H_in[966])^(data_in[199]&H_in[967])^(data_in[200]&H_in[968])^(data_in[201]&H_in[969])^(data_in[202]&H_in[970])^(data_in[203]&H_in[971])^(data_in[204]&H_in[972])^(data_in[205]&H_in[973])^(data_in[206]&H_in[974])^(data_in[207]&H_in[975])^(data_in[208]&H_in[976])^(data_in[209]&H_in[977])^(data_in[210]&H_in[978])^(data_in[211]&H_in[979])^(data_in[212]&H_in[980])^(data_in[213]&H_in[981])^(data_in[214]&H_in[982])^(data_in[215]&H_in[983])^(data_in[216]&H_in[984])^(data_in[217]&H_in[985])^(data_in[218]&H_in[986])^(data_in[219]&H_in[987])^(data_in[220]&H_in[988])^(data_in[221]&H_in[989])^(data_in[222]&H_in[990])^(data_in[223]&H_in[991])^(data_in[224]&H_in[992])^(data_in[225]&H_in[993])^(data_in[226]&H_in[994])^(data_in[227]&H_in[995])^(data_in[228]&H_in[996])^(data_in[229]&H_in[997])^(data_in[230]&H_in[998])^(data_in[231]&H_in[999])^(data_in[232]&H_in[1000])^(data_in[233]&H_in[1001])^(data_in[234]&H_in[1002])^(data_in[235]&H_in[1003])^(data_in[236]&H_in[1004])^(data_in[237]&H_in[1005])^(data_in[238]&H_in[1006])^(data_in[239]&H_in[1007])^(data_in[240]&H_in[1008])^(data_in[241]&H_in[1009])^(data_in[242]&H_in[1010])^(data_in[243]&H_in[1011])^(data_in[244]&H_in[1012])^(data_in[245]&H_in[1013])^(data_in[246]&H_in[1014])^(data_in[247]&H_in[1015])^(data_in[248]&H_in[1016])^(data_in[249]&H_in[1017])^(data_in[250]&H_in[1018])^(data_in[251]&H_in[1019])^(data_in[252]&H_in[1020])^(data_in[253]&H_in[1021])^(data_in[254]&H_in[1022])^(data_in[255]&H_in[1023]);
         data_out[4]<=(data_in[0]&H_in[1024])^(data_in[1]&H_in[1025])^(data_in[2]&H_in[1026])^(data_in[3]&H_in[1027])^(data_in[4]&H_in[1028])^(data_in[5]&H_in[1029])^(data_in[6]&H_in[1030])^(data_in[7]&H_in[1031])^(data_in[8]&H_in[1032])^(data_in[9]&H_in[1033])^(data_in[10]&H_in[1034])^(data_in[11]&H_in[1035])^(data_in[12]&H_in[1036])^(data_in[13]&H_in[1037])^(data_in[14]&H_in[1038])^(data_in[15]&H_in[1039])^(data_in[16]&H_in[1040])^(data_in[17]&H_in[1041])^(data_in[18]&H_in[1042])^(data_in[19]&H_in[1043])^(data_in[20]&H_in[1044])^(data_in[21]&H_in[1045])^(data_in[22]&H_in[1046])^(data_in[23]&H_in[1047])^(data_in[24]&H_in[1048])^(data_in[25]&H_in[1049])^(data_in[26]&H_in[1050])^(data_in[27]&H_in[1051])^(data_in[28]&H_in[1052])^(data_in[29]&H_in[1053])^(data_in[30]&H_in[1054])^(data_in[31]&H_in[1055])^(data_in[32]&H_in[1056])^(data_in[33]&H_in[1057])^(data_in[34]&H_in[1058])^(data_in[35]&H_in[1059])^(data_in[36]&H_in[1060])^(data_in[37]&H_in[1061])^(data_in[38]&H_in[1062])^(data_in[39]&H_in[1063])^(data_in[40]&H_in[1064])^(data_in[41]&H_in[1065])^(data_in[42]&H_in[1066])^(data_in[43]&H_in[1067])^(data_in[44]&H_in[1068])^(data_in[45]&H_in[1069])^(data_in[46]&H_in[1070])^(data_in[47]&H_in[1071])^(data_in[48]&H_in[1072])^(data_in[49]&H_in[1073])^(data_in[50]&H_in[1074])^(data_in[51]&H_in[1075])^(data_in[52]&H_in[1076])^(data_in[53]&H_in[1077])^(data_in[54]&H_in[1078])^(data_in[55]&H_in[1079])^(data_in[56]&H_in[1080])^(data_in[57]&H_in[1081])^(data_in[58]&H_in[1082])^(data_in[59]&H_in[1083])^(data_in[60]&H_in[1084])^(data_in[61]&H_in[1085])^(data_in[62]&H_in[1086])^(data_in[63]&H_in[1087])^(data_in[64]&H_in[1088])^(data_in[65]&H_in[1089])^(data_in[66]&H_in[1090])^(data_in[67]&H_in[1091])^(data_in[68]&H_in[1092])^(data_in[69]&H_in[1093])^(data_in[70]&H_in[1094])^(data_in[71]&H_in[1095])^(data_in[72]&H_in[1096])^(data_in[73]&H_in[1097])^(data_in[74]&H_in[1098])^(data_in[75]&H_in[1099])^(data_in[76]&H_in[1100])^(data_in[77]&H_in[1101])^(data_in[78]&H_in[1102])^(data_in[79]&H_in[1103])^(data_in[80]&H_in[1104])^(data_in[81]&H_in[1105])^(data_in[82]&H_in[1106])^(data_in[83]&H_in[1107])^(data_in[84]&H_in[1108])^(data_in[85]&H_in[1109])^(data_in[86]&H_in[1110])^(data_in[87]&H_in[1111])^(data_in[88]&H_in[1112])^(data_in[89]&H_in[1113])^(data_in[90]&H_in[1114])^(data_in[91]&H_in[1115])^(data_in[92]&H_in[1116])^(data_in[93]&H_in[1117])^(data_in[94]&H_in[1118])^(data_in[95]&H_in[1119])^(data_in[96]&H_in[1120])^(data_in[97]&H_in[1121])^(data_in[98]&H_in[1122])^(data_in[99]&H_in[1123])^(data_in[100]&H_in[1124])^(data_in[101]&H_in[1125])^(data_in[102]&H_in[1126])^(data_in[103]&H_in[1127])^(data_in[104]&H_in[1128])^(data_in[105]&H_in[1129])^(data_in[106]&H_in[1130])^(data_in[107]&H_in[1131])^(data_in[108]&H_in[1132])^(data_in[109]&H_in[1133])^(data_in[110]&H_in[1134])^(data_in[111]&H_in[1135])^(data_in[112]&H_in[1136])^(data_in[113]&H_in[1137])^(data_in[114]&H_in[1138])^(data_in[115]&H_in[1139])^(data_in[116]&H_in[1140])^(data_in[117]&H_in[1141])^(data_in[118]&H_in[1142])^(data_in[119]&H_in[1143])^(data_in[120]&H_in[1144])^(data_in[121]&H_in[1145])^(data_in[122]&H_in[1146])^(data_in[123]&H_in[1147])^(data_in[124]&H_in[1148])^(data_in[125]&H_in[1149])^(data_in[126]&H_in[1150])^(data_in[127]&H_in[1151])^(data_in[128]&H_in[1152])^(data_in[129]&H_in[1153])^(data_in[130]&H_in[1154])^(data_in[131]&H_in[1155])^(data_in[132]&H_in[1156])^(data_in[133]&H_in[1157])^(data_in[134]&H_in[1158])^(data_in[135]&H_in[1159])^(data_in[136]&H_in[1160])^(data_in[137]&H_in[1161])^(data_in[138]&H_in[1162])^(data_in[139]&H_in[1163])^(data_in[140]&H_in[1164])^(data_in[141]&H_in[1165])^(data_in[142]&H_in[1166])^(data_in[143]&H_in[1167])^(data_in[144]&H_in[1168])^(data_in[145]&H_in[1169])^(data_in[146]&H_in[1170])^(data_in[147]&H_in[1171])^(data_in[148]&H_in[1172])^(data_in[149]&H_in[1173])^(data_in[150]&H_in[1174])^(data_in[151]&H_in[1175])^(data_in[152]&H_in[1176])^(data_in[153]&H_in[1177])^(data_in[154]&H_in[1178])^(data_in[155]&H_in[1179])^(data_in[156]&H_in[1180])^(data_in[157]&H_in[1181])^(data_in[158]&H_in[1182])^(data_in[159]&H_in[1183])^(data_in[160]&H_in[1184])^(data_in[161]&H_in[1185])^(data_in[162]&H_in[1186])^(data_in[163]&H_in[1187])^(data_in[164]&H_in[1188])^(data_in[165]&H_in[1189])^(data_in[166]&H_in[1190])^(data_in[167]&H_in[1191])^(data_in[168]&H_in[1192])^(data_in[169]&H_in[1193])^(data_in[170]&H_in[1194])^(data_in[171]&H_in[1195])^(data_in[172]&H_in[1196])^(data_in[173]&H_in[1197])^(data_in[174]&H_in[1198])^(data_in[175]&H_in[1199])^(data_in[176]&H_in[1200])^(data_in[177]&H_in[1201])^(data_in[178]&H_in[1202])^(data_in[179]&H_in[1203])^(data_in[180]&H_in[1204])^(data_in[181]&H_in[1205])^(data_in[182]&H_in[1206])^(data_in[183]&H_in[1207])^(data_in[184]&H_in[1208])^(data_in[185]&H_in[1209])^(data_in[186]&H_in[1210])^(data_in[187]&H_in[1211])^(data_in[188]&H_in[1212])^(data_in[189]&H_in[1213])^(data_in[190]&H_in[1214])^(data_in[191]&H_in[1215])^(data_in[192]&H_in[1216])^(data_in[193]&H_in[1217])^(data_in[194]&H_in[1218])^(data_in[195]&H_in[1219])^(data_in[196]&H_in[1220])^(data_in[197]&H_in[1221])^(data_in[198]&H_in[1222])^(data_in[199]&H_in[1223])^(data_in[200]&H_in[1224])^(data_in[201]&H_in[1225])^(data_in[202]&H_in[1226])^(data_in[203]&H_in[1227])^(data_in[204]&H_in[1228])^(data_in[205]&H_in[1229])^(data_in[206]&H_in[1230])^(data_in[207]&H_in[1231])^(data_in[208]&H_in[1232])^(data_in[209]&H_in[1233])^(data_in[210]&H_in[1234])^(data_in[211]&H_in[1235])^(data_in[212]&H_in[1236])^(data_in[213]&H_in[1237])^(data_in[214]&H_in[1238])^(data_in[215]&H_in[1239])^(data_in[216]&H_in[1240])^(data_in[217]&H_in[1241])^(data_in[218]&H_in[1242])^(data_in[219]&H_in[1243])^(data_in[220]&H_in[1244])^(data_in[221]&H_in[1245])^(data_in[222]&H_in[1246])^(data_in[223]&H_in[1247])^(data_in[224]&H_in[1248])^(data_in[225]&H_in[1249])^(data_in[226]&H_in[1250])^(data_in[227]&H_in[1251])^(data_in[228]&H_in[1252])^(data_in[229]&H_in[1253])^(data_in[230]&H_in[1254])^(data_in[231]&H_in[1255])^(data_in[232]&H_in[1256])^(data_in[233]&H_in[1257])^(data_in[234]&H_in[1258])^(data_in[235]&H_in[1259])^(data_in[236]&H_in[1260])^(data_in[237]&H_in[1261])^(data_in[238]&H_in[1262])^(data_in[239]&H_in[1263])^(data_in[240]&H_in[1264])^(data_in[241]&H_in[1265])^(data_in[242]&H_in[1266])^(data_in[243]&H_in[1267])^(data_in[244]&H_in[1268])^(data_in[245]&H_in[1269])^(data_in[246]&H_in[1270])^(data_in[247]&H_in[1271])^(data_in[248]&H_in[1272])^(data_in[249]&H_in[1273])^(data_in[250]&H_in[1274])^(data_in[251]&H_in[1275])^(data_in[252]&H_in[1276])^(data_in[253]&H_in[1277])^(data_in[254]&H_in[1278])^(data_in[255]&H_in[1279]);
         data_out[5]<=(data_in[0]&H_in[1280])^(data_in[1]&H_in[1281])^(data_in[2]&H_in[1282])^(data_in[3]&H_in[1283])^(data_in[4]&H_in[1284])^(data_in[5]&H_in[1285])^(data_in[6]&H_in[1286])^(data_in[7]&H_in[1287])^(data_in[8]&H_in[1288])^(data_in[9]&H_in[1289])^(data_in[10]&H_in[1290])^(data_in[11]&H_in[1291])^(data_in[12]&H_in[1292])^(data_in[13]&H_in[1293])^(data_in[14]&H_in[1294])^(data_in[15]&H_in[1295])^(data_in[16]&H_in[1296])^(data_in[17]&H_in[1297])^(data_in[18]&H_in[1298])^(data_in[19]&H_in[1299])^(data_in[20]&H_in[1300])^(data_in[21]&H_in[1301])^(data_in[22]&H_in[1302])^(data_in[23]&H_in[1303])^(data_in[24]&H_in[1304])^(data_in[25]&H_in[1305])^(data_in[26]&H_in[1306])^(data_in[27]&H_in[1307])^(data_in[28]&H_in[1308])^(data_in[29]&H_in[1309])^(data_in[30]&H_in[1310])^(data_in[31]&H_in[1311])^(data_in[32]&H_in[1312])^(data_in[33]&H_in[1313])^(data_in[34]&H_in[1314])^(data_in[35]&H_in[1315])^(data_in[36]&H_in[1316])^(data_in[37]&H_in[1317])^(data_in[38]&H_in[1318])^(data_in[39]&H_in[1319])^(data_in[40]&H_in[1320])^(data_in[41]&H_in[1321])^(data_in[42]&H_in[1322])^(data_in[43]&H_in[1323])^(data_in[44]&H_in[1324])^(data_in[45]&H_in[1325])^(data_in[46]&H_in[1326])^(data_in[47]&H_in[1327])^(data_in[48]&H_in[1328])^(data_in[49]&H_in[1329])^(data_in[50]&H_in[1330])^(data_in[51]&H_in[1331])^(data_in[52]&H_in[1332])^(data_in[53]&H_in[1333])^(data_in[54]&H_in[1334])^(data_in[55]&H_in[1335])^(data_in[56]&H_in[1336])^(data_in[57]&H_in[1337])^(data_in[58]&H_in[1338])^(data_in[59]&H_in[1339])^(data_in[60]&H_in[1340])^(data_in[61]&H_in[1341])^(data_in[62]&H_in[1342])^(data_in[63]&H_in[1343])^(data_in[64]&H_in[1344])^(data_in[65]&H_in[1345])^(data_in[66]&H_in[1346])^(data_in[67]&H_in[1347])^(data_in[68]&H_in[1348])^(data_in[69]&H_in[1349])^(data_in[70]&H_in[1350])^(data_in[71]&H_in[1351])^(data_in[72]&H_in[1352])^(data_in[73]&H_in[1353])^(data_in[74]&H_in[1354])^(data_in[75]&H_in[1355])^(data_in[76]&H_in[1356])^(data_in[77]&H_in[1357])^(data_in[78]&H_in[1358])^(data_in[79]&H_in[1359])^(data_in[80]&H_in[1360])^(data_in[81]&H_in[1361])^(data_in[82]&H_in[1362])^(data_in[83]&H_in[1363])^(data_in[84]&H_in[1364])^(data_in[85]&H_in[1365])^(data_in[86]&H_in[1366])^(data_in[87]&H_in[1367])^(data_in[88]&H_in[1368])^(data_in[89]&H_in[1369])^(data_in[90]&H_in[1370])^(data_in[91]&H_in[1371])^(data_in[92]&H_in[1372])^(data_in[93]&H_in[1373])^(data_in[94]&H_in[1374])^(data_in[95]&H_in[1375])^(data_in[96]&H_in[1376])^(data_in[97]&H_in[1377])^(data_in[98]&H_in[1378])^(data_in[99]&H_in[1379])^(data_in[100]&H_in[1380])^(data_in[101]&H_in[1381])^(data_in[102]&H_in[1382])^(data_in[103]&H_in[1383])^(data_in[104]&H_in[1384])^(data_in[105]&H_in[1385])^(data_in[106]&H_in[1386])^(data_in[107]&H_in[1387])^(data_in[108]&H_in[1388])^(data_in[109]&H_in[1389])^(data_in[110]&H_in[1390])^(data_in[111]&H_in[1391])^(data_in[112]&H_in[1392])^(data_in[113]&H_in[1393])^(data_in[114]&H_in[1394])^(data_in[115]&H_in[1395])^(data_in[116]&H_in[1396])^(data_in[117]&H_in[1397])^(data_in[118]&H_in[1398])^(data_in[119]&H_in[1399])^(data_in[120]&H_in[1400])^(data_in[121]&H_in[1401])^(data_in[122]&H_in[1402])^(data_in[123]&H_in[1403])^(data_in[124]&H_in[1404])^(data_in[125]&H_in[1405])^(data_in[126]&H_in[1406])^(data_in[127]&H_in[1407])^(data_in[128]&H_in[1408])^(data_in[129]&H_in[1409])^(data_in[130]&H_in[1410])^(data_in[131]&H_in[1411])^(data_in[132]&H_in[1412])^(data_in[133]&H_in[1413])^(data_in[134]&H_in[1414])^(data_in[135]&H_in[1415])^(data_in[136]&H_in[1416])^(data_in[137]&H_in[1417])^(data_in[138]&H_in[1418])^(data_in[139]&H_in[1419])^(data_in[140]&H_in[1420])^(data_in[141]&H_in[1421])^(data_in[142]&H_in[1422])^(data_in[143]&H_in[1423])^(data_in[144]&H_in[1424])^(data_in[145]&H_in[1425])^(data_in[146]&H_in[1426])^(data_in[147]&H_in[1427])^(data_in[148]&H_in[1428])^(data_in[149]&H_in[1429])^(data_in[150]&H_in[1430])^(data_in[151]&H_in[1431])^(data_in[152]&H_in[1432])^(data_in[153]&H_in[1433])^(data_in[154]&H_in[1434])^(data_in[155]&H_in[1435])^(data_in[156]&H_in[1436])^(data_in[157]&H_in[1437])^(data_in[158]&H_in[1438])^(data_in[159]&H_in[1439])^(data_in[160]&H_in[1440])^(data_in[161]&H_in[1441])^(data_in[162]&H_in[1442])^(data_in[163]&H_in[1443])^(data_in[164]&H_in[1444])^(data_in[165]&H_in[1445])^(data_in[166]&H_in[1446])^(data_in[167]&H_in[1447])^(data_in[168]&H_in[1448])^(data_in[169]&H_in[1449])^(data_in[170]&H_in[1450])^(data_in[171]&H_in[1451])^(data_in[172]&H_in[1452])^(data_in[173]&H_in[1453])^(data_in[174]&H_in[1454])^(data_in[175]&H_in[1455])^(data_in[176]&H_in[1456])^(data_in[177]&H_in[1457])^(data_in[178]&H_in[1458])^(data_in[179]&H_in[1459])^(data_in[180]&H_in[1460])^(data_in[181]&H_in[1461])^(data_in[182]&H_in[1462])^(data_in[183]&H_in[1463])^(data_in[184]&H_in[1464])^(data_in[185]&H_in[1465])^(data_in[186]&H_in[1466])^(data_in[187]&H_in[1467])^(data_in[188]&H_in[1468])^(data_in[189]&H_in[1469])^(data_in[190]&H_in[1470])^(data_in[191]&H_in[1471])^(data_in[192]&H_in[1472])^(data_in[193]&H_in[1473])^(data_in[194]&H_in[1474])^(data_in[195]&H_in[1475])^(data_in[196]&H_in[1476])^(data_in[197]&H_in[1477])^(data_in[198]&H_in[1478])^(data_in[199]&H_in[1479])^(data_in[200]&H_in[1480])^(data_in[201]&H_in[1481])^(data_in[202]&H_in[1482])^(data_in[203]&H_in[1483])^(data_in[204]&H_in[1484])^(data_in[205]&H_in[1485])^(data_in[206]&H_in[1486])^(data_in[207]&H_in[1487])^(data_in[208]&H_in[1488])^(data_in[209]&H_in[1489])^(data_in[210]&H_in[1490])^(data_in[211]&H_in[1491])^(data_in[212]&H_in[1492])^(data_in[213]&H_in[1493])^(data_in[214]&H_in[1494])^(data_in[215]&H_in[1495])^(data_in[216]&H_in[1496])^(data_in[217]&H_in[1497])^(data_in[218]&H_in[1498])^(data_in[219]&H_in[1499])^(data_in[220]&H_in[1500])^(data_in[221]&H_in[1501])^(data_in[222]&H_in[1502])^(data_in[223]&H_in[1503])^(data_in[224]&H_in[1504])^(data_in[225]&H_in[1505])^(data_in[226]&H_in[1506])^(data_in[227]&H_in[1507])^(data_in[228]&H_in[1508])^(data_in[229]&H_in[1509])^(data_in[230]&H_in[1510])^(data_in[231]&H_in[1511])^(data_in[232]&H_in[1512])^(data_in[233]&H_in[1513])^(data_in[234]&H_in[1514])^(data_in[235]&H_in[1515])^(data_in[236]&H_in[1516])^(data_in[237]&H_in[1517])^(data_in[238]&H_in[1518])^(data_in[239]&H_in[1519])^(data_in[240]&H_in[1520])^(data_in[241]&H_in[1521])^(data_in[242]&H_in[1522])^(data_in[243]&H_in[1523])^(data_in[244]&H_in[1524])^(data_in[245]&H_in[1525])^(data_in[246]&H_in[1526])^(data_in[247]&H_in[1527])^(data_in[248]&H_in[1528])^(data_in[249]&H_in[1529])^(data_in[250]&H_in[1530])^(data_in[251]&H_in[1531])^(data_in[252]&H_in[1532])^(data_in[253]&H_in[1533])^(data_in[254]&H_in[1534])^(data_in[255]&H_in[1535]);
         data_out[6]<=(data_in[0]&H_in[1536])^(data_in[1]&H_in[1537])^(data_in[2]&H_in[1538])^(data_in[3]&H_in[1539])^(data_in[4]&H_in[1540])^(data_in[5]&H_in[1541])^(data_in[6]&H_in[1542])^(data_in[7]&H_in[1543])^(data_in[8]&H_in[1544])^(data_in[9]&H_in[1545])^(data_in[10]&H_in[1546])^(data_in[11]&H_in[1547])^(data_in[12]&H_in[1548])^(data_in[13]&H_in[1549])^(data_in[14]&H_in[1550])^(data_in[15]&H_in[1551])^(data_in[16]&H_in[1552])^(data_in[17]&H_in[1553])^(data_in[18]&H_in[1554])^(data_in[19]&H_in[1555])^(data_in[20]&H_in[1556])^(data_in[21]&H_in[1557])^(data_in[22]&H_in[1558])^(data_in[23]&H_in[1559])^(data_in[24]&H_in[1560])^(data_in[25]&H_in[1561])^(data_in[26]&H_in[1562])^(data_in[27]&H_in[1563])^(data_in[28]&H_in[1564])^(data_in[29]&H_in[1565])^(data_in[30]&H_in[1566])^(data_in[31]&H_in[1567])^(data_in[32]&H_in[1568])^(data_in[33]&H_in[1569])^(data_in[34]&H_in[1570])^(data_in[35]&H_in[1571])^(data_in[36]&H_in[1572])^(data_in[37]&H_in[1573])^(data_in[38]&H_in[1574])^(data_in[39]&H_in[1575])^(data_in[40]&H_in[1576])^(data_in[41]&H_in[1577])^(data_in[42]&H_in[1578])^(data_in[43]&H_in[1579])^(data_in[44]&H_in[1580])^(data_in[45]&H_in[1581])^(data_in[46]&H_in[1582])^(data_in[47]&H_in[1583])^(data_in[48]&H_in[1584])^(data_in[49]&H_in[1585])^(data_in[50]&H_in[1586])^(data_in[51]&H_in[1587])^(data_in[52]&H_in[1588])^(data_in[53]&H_in[1589])^(data_in[54]&H_in[1590])^(data_in[55]&H_in[1591])^(data_in[56]&H_in[1592])^(data_in[57]&H_in[1593])^(data_in[58]&H_in[1594])^(data_in[59]&H_in[1595])^(data_in[60]&H_in[1596])^(data_in[61]&H_in[1597])^(data_in[62]&H_in[1598])^(data_in[63]&H_in[1599])^(data_in[64]&H_in[1600])^(data_in[65]&H_in[1601])^(data_in[66]&H_in[1602])^(data_in[67]&H_in[1603])^(data_in[68]&H_in[1604])^(data_in[69]&H_in[1605])^(data_in[70]&H_in[1606])^(data_in[71]&H_in[1607])^(data_in[72]&H_in[1608])^(data_in[73]&H_in[1609])^(data_in[74]&H_in[1610])^(data_in[75]&H_in[1611])^(data_in[76]&H_in[1612])^(data_in[77]&H_in[1613])^(data_in[78]&H_in[1614])^(data_in[79]&H_in[1615])^(data_in[80]&H_in[1616])^(data_in[81]&H_in[1617])^(data_in[82]&H_in[1618])^(data_in[83]&H_in[1619])^(data_in[84]&H_in[1620])^(data_in[85]&H_in[1621])^(data_in[86]&H_in[1622])^(data_in[87]&H_in[1623])^(data_in[88]&H_in[1624])^(data_in[89]&H_in[1625])^(data_in[90]&H_in[1626])^(data_in[91]&H_in[1627])^(data_in[92]&H_in[1628])^(data_in[93]&H_in[1629])^(data_in[94]&H_in[1630])^(data_in[95]&H_in[1631])^(data_in[96]&H_in[1632])^(data_in[97]&H_in[1633])^(data_in[98]&H_in[1634])^(data_in[99]&H_in[1635])^(data_in[100]&H_in[1636])^(data_in[101]&H_in[1637])^(data_in[102]&H_in[1638])^(data_in[103]&H_in[1639])^(data_in[104]&H_in[1640])^(data_in[105]&H_in[1641])^(data_in[106]&H_in[1642])^(data_in[107]&H_in[1643])^(data_in[108]&H_in[1644])^(data_in[109]&H_in[1645])^(data_in[110]&H_in[1646])^(data_in[111]&H_in[1647])^(data_in[112]&H_in[1648])^(data_in[113]&H_in[1649])^(data_in[114]&H_in[1650])^(data_in[115]&H_in[1651])^(data_in[116]&H_in[1652])^(data_in[117]&H_in[1653])^(data_in[118]&H_in[1654])^(data_in[119]&H_in[1655])^(data_in[120]&H_in[1656])^(data_in[121]&H_in[1657])^(data_in[122]&H_in[1658])^(data_in[123]&H_in[1659])^(data_in[124]&H_in[1660])^(data_in[125]&H_in[1661])^(data_in[126]&H_in[1662])^(data_in[127]&H_in[1663])^(data_in[128]&H_in[1664])^(data_in[129]&H_in[1665])^(data_in[130]&H_in[1666])^(data_in[131]&H_in[1667])^(data_in[132]&H_in[1668])^(data_in[133]&H_in[1669])^(data_in[134]&H_in[1670])^(data_in[135]&H_in[1671])^(data_in[136]&H_in[1672])^(data_in[137]&H_in[1673])^(data_in[138]&H_in[1674])^(data_in[139]&H_in[1675])^(data_in[140]&H_in[1676])^(data_in[141]&H_in[1677])^(data_in[142]&H_in[1678])^(data_in[143]&H_in[1679])^(data_in[144]&H_in[1680])^(data_in[145]&H_in[1681])^(data_in[146]&H_in[1682])^(data_in[147]&H_in[1683])^(data_in[148]&H_in[1684])^(data_in[149]&H_in[1685])^(data_in[150]&H_in[1686])^(data_in[151]&H_in[1687])^(data_in[152]&H_in[1688])^(data_in[153]&H_in[1689])^(data_in[154]&H_in[1690])^(data_in[155]&H_in[1691])^(data_in[156]&H_in[1692])^(data_in[157]&H_in[1693])^(data_in[158]&H_in[1694])^(data_in[159]&H_in[1695])^(data_in[160]&H_in[1696])^(data_in[161]&H_in[1697])^(data_in[162]&H_in[1698])^(data_in[163]&H_in[1699])^(data_in[164]&H_in[1700])^(data_in[165]&H_in[1701])^(data_in[166]&H_in[1702])^(data_in[167]&H_in[1703])^(data_in[168]&H_in[1704])^(data_in[169]&H_in[1705])^(data_in[170]&H_in[1706])^(data_in[171]&H_in[1707])^(data_in[172]&H_in[1708])^(data_in[173]&H_in[1709])^(data_in[174]&H_in[1710])^(data_in[175]&H_in[1711])^(data_in[176]&H_in[1712])^(data_in[177]&H_in[1713])^(data_in[178]&H_in[1714])^(data_in[179]&H_in[1715])^(data_in[180]&H_in[1716])^(data_in[181]&H_in[1717])^(data_in[182]&H_in[1718])^(data_in[183]&H_in[1719])^(data_in[184]&H_in[1720])^(data_in[185]&H_in[1721])^(data_in[186]&H_in[1722])^(data_in[187]&H_in[1723])^(data_in[188]&H_in[1724])^(data_in[189]&H_in[1725])^(data_in[190]&H_in[1726])^(data_in[191]&H_in[1727])^(data_in[192]&H_in[1728])^(data_in[193]&H_in[1729])^(data_in[194]&H_in[1730])^(data_in[195]&H_in[1731])^(data_in[196]&H_in[1732])^(data_in[197]&H_in[1733])^(data_in[198]&H_in[1734])^(data_in[199]&H_in[1735])^(data_in[200]&H_in[1736])^(data_in[201]&H_in[1737])^(data_in[202]&H_in[1738])^(data_in[203]&H_in[1739])^(data_in[204]&H_in[1740])^(data_in[205]&H_in[1741])^(data_in[206]&H_in[1742])^(data_in[207]&H_in[1743])^(data_in[208]&H_in[1744])^(data_in[209]&H_in[1745])^(data_in[210]&H_in[1746])^(data_in[211]&H_in[1747])^(data_in[212]&H_in[1748])^(data_in[213]&H_in[1749])^(data_in[214]&H_in[1750])^(data_in[215]&H_in[1751])^(data_in[216]&H_in[1752])^(data_in[217]&H_in[1753])^(data_in[218]&H_in[1754])^(data_in[219]&H_in[1755])^(data_in[220]&H_in[1756])^(data_in[221]&H_in[1757])^(data_in[222]&H_in[1758])^(data_in[223]&H_in[1759])^(data_in[224]&H_in[1760])^(data_in[225]&H_in[1761])^(data_in[226]&H_in[1762])^(data_in[227]&H_in[1763])^(data_in[228]&H_in[1764])^(data_in[229]&H_in[1765])^(data_in[230]&H_in[1766])^(data_in[231]&H_in[1767])^(data_in[232]&H_in[1768])^(data_in[233]&H_in[1769])^(data_in[234]&H_in[1770])^(data_in[235]&H_in[1771])^(data_in[236]&H_in[1772])^(data_in[237]&H_in[1773])^(data_in[238]&H_in[1774])^(data_in[239]&H_in[1775])^(data_in[240]&H_in[1776])^(data_in[241]&H_in[1777])^(data_in[242]&H_in[1778])^(data_in[243]&H_in[1779])^(data_in[244]&H_in[1780])^(data_in[245]&H_in[1781])^(data_in[246]&H_in[1782])^(data_in[247]&H_in[1783])^(data_in[248]&H_in[1784])^(data_in[249]&H_in[1785])^(data_in[250]&H_in[1786])^(data_in[251]&H_in[1787])^(data_in[252]&H_in[1788])^(data_in[253]&H_in[1789])^(data_in[254]&H_in[1790])^(data_in[255]&H_in[1791]);
         data_out[7]<=(data_in[0]&H_in[1792])^(data_in[1]&H_in[1793])^(data_in[2]&H_in[1794])^(data_in[3]&H_in[1795])^(data_in[4]&H_in[1796])^(data_in[5]&H_in[1797])^(data_in[6]&H_in[1798])^(data_in[7]&H_in[1799])^(data_in[8]&H_in[1800])^(data_in[9]&H_in[1801])^(data_in[10]&H_in[1802])^(data_in[11]&H_in[1803])^(data_in[12]&H_in[1804])^(data_in[13]&H_in[1805])^(data_in[14]&H_in[1806])^(data_in[15]&H_in[1807])^(data_in[16]&H_in[1808])^(data_in[17]&H_in[1809])^(data_in[18]&H_in[1810])^(data_in[19]&H_in[1811])^(data_in[20]&H_in[1812])^(data_in[21]&H_in[1813])^(data_in[22]&H_in[1814])^(data_in[23]&H_in[1815])^(data_in[24]&H_in[1816])^(data_in[25]&H_in[1817])^(data_in[26]&H_in[1818])^(data_in[27]&H_in[1819])^(data_in[28]&H_in[1820])^(data_in[29]&H_in[1821])^(data_in[30]&H_in[1822])^(data_in[31]&H_in[1823])^(data_in[32]&H_in[1824])^(data_in[33]&H_in[1825])^(data_in[34]&H_in[1826])^(data_in[35]&H_in[1827])^(data_in[36]&H_in[1828])^(data_in[37]&H_in[1829])^(data_in[38]&H_in[1830])^(data_in[39]&H_in[1831])^(data_in[40]&H_in[1832])^(data_in[41]&H_in[1833])^(data_in[42]&H_in[1834])^(data_in[43]&H_in[1835])^(data_in[44]&H_in[1836])^(data_in[45]&H_in[1837])^(data_in[46]&H_in[1838])^(data_in[47]&H_in[1839])^(data_in[48]&H_in[1840])^(data_in[49]&H_in[1841])^(data_in[50]&H_in[1842])^(data_in[51]&H_in[1843])^(data_in[52]&H_in[1844])^(data_in[53]&H_in[1845])^(data_in[54]&H_in[1846])^(data_in[55]&H_in[1847])^(data_in[56]&H_in[1848])^(data_in[57]&H_in[1849])^(data_in[58]&H_in[1850])^(data_in[59]&H_in[1851])^(data_in[60]&H_in[1852])^(data_in[61]&H_in[1853])^(data_in[62]&H_in[1854])^(data_in[63]&H_in[1855])^(data_in[64]&H_in[1856])^(data_in[65]&H_in[1857])^(data_in[66]&H_in[1858])^(data_in[67]&H_in[1859])^(data_in[68]&H_in[1860])^(data_in[69]&H_in[1861])^(data_in[70]&H_in[1862])^(data_in[71]&H_in[1863])^(data_in[72]&H_in[1864])^(data_in[73]&H_in[1865])^(data_in[74]&H_in[1866])^(data_in[75]&H_in[1867])^(data_in[76]&H_in[1868])^(data_in[77]&H_in[1869])^(data_in[78]&H_in[1870])^(data_in[79]&H_in[1871])^(data_in[80]&H_in[1872])^(data_in[81]&H_in[1873])^(data_in[82]&H_in[1874])^(data_in[83]&H_in[1875])^(data_in[84]&H_in[1876])^(data_in[85]&H_in[1877])^(data_in[86]&H_in[1878])^(data_in[87]&H_in[1879])^(data_in[88]&H_in[1880])^(data_in[89]&H_in[1881])^(data_in[90]&H_in[1882])^(data_in[91]&H_in[1883])^(data_in[92]&H_in[1884])^(data_in[93]&H_in[1885])^(data_in[94]&H_in[1886])^(data_in[95]&H_in[1887])^(data_in[96]&H_in[1888])^(data_in[97]&H_in[1889])^(data_in[98]&H_in[1890])^(data_in[99]&H_in[1891])^(data_in[100]&H_in[1892])^(data_in[101]&H_in[1893])^(data_in[102]&H_in[1894])^(data_in[103]&H_in[1895])^(data_in[104]&H_in[1896])^(data_in[105]&H_in[1897])^(data_in[106]&H_in[1898])^(data_in[107]&H_in[1899])^(data_in[108]&H_in[1900])^(data_in[109]&H_in[1901])^(data_in[110]&H_in[1902])^(data_in[111]&H_in[1903])^(data_in[112]&H_in[1904])^(data_in[113]&H_in[1905])^(data_in[114]&H_in[1906])^(data_in[115]&H_in[1907])^(data_in[116]&H_in[1908])^(data_in[117]&H_in[1909])^(data_in[118]&H_in[1910])^(data_in[119]&H_in[1911])^(data_in[120]&H_in[1912])^(data_in[121]&H_in[1913])^(data_in[122]&H_in[1914])^(data_in[123]&H_in[1915])^(data_in[124]&H_in[1916])^(data_in[125]&H_in[1917])^(data_in[126]&H_in[1918])^(data_in[127]&H_in[1919])^(data_in[128]&H_in[1920])^(data_in[129]&H_in[1921])^(data_in[130]&H_in[1922])^(data_in[131]&H_in[1923])^(data_in[132]&H_in[1924])^(data_in[133]&H_in[1925])^(data_in[134]&H_in[1926])^(data_in[135]&H_in[1927])^(data_in[136]&H_in[1928])^(data_in[137]&H_in[1929])^(data_in[138]&H_in[1930])^(data_in[139]&H_in[1931])^(data_in[140]&H_in[1932])^(data_in[141]&H_in[1933])^(data_in[142]&H_in[1934])^(data_in[143]&H_in[1935])^(data_in[144]&H_in[1936])^(data_in[145]&H_in[1937])^(data_in[146]&H_in[1938])^(data_in[147]&H_in[1939])^(data_in[148]&H_in[1940])^(data_in[149]&H_in[1941])^(data_in[150]&H_in[1942])^(data_in[151]&H_in[1943])^(data_in[152]&H_in[1944])^(data_in[153]&H_in[1945])^(data_in[154]&H_in[1946])^(data_in[155]&H_in[1947])^(data_in[156]&H_in[1948])^(data_in[157]&H_in[1949])^(data_in[158]&H_in[1950])^(data_in[159]&H_in[1951])^(data_in[160]&H_in[1952])^(data_in[161]&H_in[1953])^(data_in[162]&H_in[1954])^(data_in[163]&H_in[1955])^(data_in[164]&H_in[1956])^(data_in[165]&H_in[1957])^(data_in[166]&H_in[1958])^(data_in[167]&H_in[1959])^(data_in[168]&H_in[1960])^(data_in[169]&H_in[1961])^(data_in[170]&H_in[1962])^(data_in[171]&H_in[1963])^(data_in[172]&H_in[1964])^(data_in[173]&H_in[1965])^(data_in[174]&H_in[1966])^(data_in[175]&H_in[1967])^(data_in[176]&H_in[1968])^(data_in[177]&H_in[1969])^(data_in[178]&H_in[1970])^(data_in[179]&H_in[1971])^(data_in[180]&H_in[1972])^(data_in[181]&H_in[1973])^(data_in[182]&H_in[1974])^(data_in[183]&H_in[1975])^(data_in[184]&H_in[1976])^(data_in[185]&H_in[1977])^(data_in[186]&H_in[1978])^(data_in[187]&H_in[1979])^(data_in[188]&H_in[1980])^(data_in[189]&H_in[1981])^(data_in[190]&H_in[1982])^(data_in[191]&H_in[1983])^(data_in[192]&H_in[1984])^(data_in[193]&H_in[1985])^(data_in[194]&H_in[1986])^(data_in[195]&H_in[1987])^(data_in[196]&H_in[1988])^(data_in[197]&H_in[1989])^(data_in[198]&H_in[1990])^(data_in[199]&H_in[1991])^(data_in[200]&H_in[1992])^(data_in[201]&H_in[1993])^(data_in[202]&H_in[1994])^(data_in[203]&H_in[1995])^(data_in[204]&H_in[1996])^(data_in[205]&H_in[1997])^(data_in[206]&H_in[1998])^(data_in[207]&H_in[1999])^(data_in[208]&H_in[2000])^(data_in[209]&H_in[2001])^(data_in[210]&H_in[2002])^(data_in[211]&H_in[2003])^(data_in[212]&H_in[2004])^(data_in[213]&H_in[2005])^(data_in[214]&H_in[2006])^(data_in[215]&H_in[2007])^(data_in[216]&H_in[2008])^(data_in[217]&H_in[2009])^(data_in[218]&H_in[2010])^(data_in[219]&H_in[2011])^(data_in[220]&H_in[2012])^(data_in[221]&H_in[2013])^(data_in[222]&H_in[2014])^(data_in[223]&H_in[2015])^(data_in[224]&H_in[2016])^(data_in[225]&H_in[2017])^(data_in[226]&H_in[2018])^(data_in[227]&H_in[2019])^(data_in[228]&H_in[2020])^(data_in[229]&H_in[2021])^(data_in[230]&H_in[2022])^(data_in[231]&H_in[2023])^(data_in[232]&H_in[2024])^(data_in[233]&H_in[2025])^(data_in[234]&H_in[2026])^(data_in[235]&H_in[2027])^(data_in[236]&H_in[2028])^(data_in[237]&H_in[2029])^(data_in[238]&H_in[2030])^(data_in[239]&H_in[2031])^(data_in[240]&H_in[2032])^(data_in[241]&H_in[2033])^(data_in[242]&H_in[2034])^(data_in[243]&H_in[2035])^(data_in[244]&H_in[2036])^(data_in[245]&H_in[2037])^(data_in[246]&H_in[2038])^(data_in[247]&H_in[2039])^(data_in[248]&H_in[2040])^(data_in[249]&H_in[2041])^(data_in[250]&H_in[2042])^(data_in[251]&H_in[2043])^(data_in[252]&H_in[2044])^(data_in[253]&H_in[2045])^(data_in[254]&H_in[2046])^(data_in[255]&H_in[2047]);
         data_out[8]<=(data_in[0]&H_in[2048])^(data_in[1]&H_in[2049])^(data_in[2]&H_in[2050])^(data_in[3]&H_in[2051])^(data_in[4]&H_in[2052])^(data_in[5]&H_in[2053])^(data_in[6]&H_in[2054])^(data_in[7]&H_in[2055])^(data_in[8]&H_in[2056])^(data_in[9]&H_in[2057])^(data_in[10]&H_in[2058])^(data_in[11]&H_in[2059])^(data_in[12]&H_in[2060])^(data_in[13]&H_in[2061])^(data_in[14]&H_in[2062])^(data_in[15]&H_in[2063])^(data_in[16]&H_in[2064])^(data_in[17]&H_in[2065])^(data_in[18]&H_in[2066])^(data_in[19]&H_in[2067])^(data_in[20]&H_in[2068])^(data_in[21]&H_in[2069])^(data_in[22]&H_in[2070])^(data_in[23]&H_in[2071])^(data_in[24]&H_in[2072])^(data_in[25]&H_in[2073])^(data_in[26]&H_in[2074])^(data_in[27]&H_in[2075])^(data_in[28]&H_in[2076])^(data_in[29]&H_in[2077])^(data_in[30]&H_in[2078])^(data_in[31]&H_in[2079])^(data_in[32]&H_in[2080])^(data_in[33]&H_in[2081])^(data_in[34]&H_in[2082])^(data_in[35]&H_in[2083])^(data_in[36]&H_in[2084])^(data_in[37]&H_in[2085])^(data_in[38]&H_in[2086])^(data_in[39]&H_in[2087])^(data_in[40]&H_in[2088])^(data_in[41]&H_in[2089])^(data_in[42]&H_in[2090])^(data_in[43]&H_in[2091])^(data_in[44]&H_in[2092])^(data_in[45]&H_in[2093])^(data_in[46]&H_in[2094])^(data_in[47]&H_in[2095])^(data_in[48]&H_in[2096])^(data_in[49]&H_in[2097])^(data_in[50]&H_in[2098])^(data_in[51]&H_in[2099])^(data_in[52]&H_in[2100])^(data_in[53]&H_in[2101])^(data_in[54]&H_in[2102])^(data_in[55]&H_in[2103])^(data_in[56]&H_in[2104])^(data_in[57]&H_in[2105])^(data_in[58]&H_in[2106])^(data_in[59]&H_in[2107])^(data_in[60]&H_in[2108])^(data_in[61]&H_in[2109])^(data_in[62]&H_in[2110])^(data_in[63]&H_in[2111])^(data_in[64]&H_in[2112])^(data_in[65]&H_in[2113])^(data_in[66]&H_in[2114])^(data_in[67]&H_in[2115])^(data_in[68]&H_in[2116])^(data_in[69]&H_in[2117])^(data_in[70]&H_in[2118])^(data_in[71]&H_in[2119])^(data_in[72]&H_in[2120])^(data_in[73]&H_in[2121])^(data_in[74]&H_in[2122])^(data_in[75]&H_in[2123])^(data_in[76]&H_in[2124])^(data_in[77]&H_in[2125])^(data_in[78]&H_in[2126])^(data_in[79]&H_in[2127])^(data_in[80]&H_in[2128])^(data_in[81]&H_in[2129])^(data_in[82]&H_in[2130])^(data_in[83]&H_in[2131])^(data_in[84]&H_in[2132])^(data_in[85]&H_in[2133])^(data_in[86]&H_in[2134])^(data_in[87]&H_in[2135])^(data_in[88]&H_in[2136])^(data_in[89]&H_in[2137])^(data_in[90]&H_in[2138])^(data_in[91]&H_in[2139])^(data_in[92]&H_in[2140])^(data_in[93]&H_in[2141])^(data_in[94]&H_in[2142])^(data_in[95]&H_in[2143])^(data_in[96]&H_in[2144])^(data_in[97]&H_in[2145])^(data_in[98]&H_in[2146])^(data_in[99]&H_in[2147])^(data_in[100]&H_in[2148])^(data_in[101]&H_in[2149])^(data_in[102]&H_in[2150])^(data_in[103]&H_in[2151])^(data_in[104]&H_in[2152])^(data_in[105]&H_in[2153])^(data_in[106]&H_in[2154])^(data_in[107]&H_in[2155])^(data_in[108]&H_in[2156])^(data_in[109]&H_in[2157])^(data_in[110]&H_in[2158])^(data_in[111]&H_in[2159])^(data_in[112]&H_in[2160])^(data_in[113]&H_in[2161])^(data_in[114]&H_in[2162])^(data_in[115]&H_in[2163])^(data_in[116]&H_in[2164])^(data_in[117]&H_in[2165])^(data_in[118]&H_in[2166])^(data_in[119]&H_in[2167])^(data_in[120]&H_in[2168])^(data_in[121]&H_in[2169])^(data_in[122]&H_in[2170])^(data_in[123]&H_in[2171])^(data_in[124]&H_in[2172])^(data_in[125]&H_in[2173])^(data_in[126]&H_in[2174])^(data_in[127]&H_in[2175])^(data_in[128]&H_in[2176])^(data_in[129]&H_in[2177])^(data_in[130]&H_in[2178])^(data_in[131]&H_in[2179])^(data_in[132]&H_in[2180])^(data_in[133]&H_in[2181])^(data_in[134]&H_in[2182])^(data_in[135]&H_in[2183])^(data_in[136]&H_in[2184])^(data_in[137]&H_in[2185])^(data_in[138]&H_in[2186])^(data_in[139]&H_in[2187])^(data_in[140]&H_in[2188])^(data_in[141]&H_in[2189])^(data_in[142]&H_in[2190])^(data_in[143]&H_in[2191])^(data_in[144]&H_in[2192])^(data_in[145]&H_in[2193])^(data_in[146]&H_in[2194])^(data_in[147]&H_in[2195])^(data_in[148]&H_in[2196])^(data_in[149]&H_in[2197])^(data_in[150]&H_in[2198])^(data_in[151]&H_in[2199])^(data_in[152]&H_in[2200])^(data_in[153]&H_in[2201])^(data_in[154]&H_in[2202])^(data_in[155]&H_in[2203])^(data_in[156]&H_in[2204])^(data_in[157]&H_in[2205])^(data_in[158]&H_in[2206])^(data_in[159]&H_in[2207])^(data_in[160]&H_in[2208])^(data_in[161]&H_in[2209])^(data_in[162]&H_in[2210])^(data_in[163]&H_in[2211])^(data_in[164]&H_in[2212])^(data_in[165]&H_in[2213])^(data_in[166]&H_in[2214])^(data_in[167]&H_in[2215])^(data_in[168]&H_in[2216])^(data_in[169]&H_in[2217])^(data_in[170]&H_in[2218])^(data_in[171]&H_in[2219])^(data_in[172]&H_in[2220])^(data_in[173]&H_in[2221])^(data_in[174]&H_in[2222])^(data_in[175]&H_in[2223])^(data_in[176]&H_in[2224])^(data_in[177]&H_in[2225])^(data_in[178]&H_in[2226])^(data_in[179]&H_in[2227])^(data_in[180]&H_in[2228])^(data_in[181]&H_in[2229])^(data_in[182]&H_in[2230])^(data_in[183]&H_in[2231])^(data_in[184]&H_in[2232])^(data_in[185]&H_in[2233])^(data_in[186]&H_in[2234])^(data_in[187]&H_in[2235])^(data_in[188]&H_in[2236])^(data_in[189]&H_in[2237])^(data_in[190]&H_in[2238])^(data_in[191]&H_in[2239])^(data_in[192]&H_in[2240])^(data_in[193]&H_in[2241])^(data_in[194]&H_in[2242])^(data_in[195]&H_in[2243])^(data_in[196]&H_in[2244])^(data_in[197]&H_in[2245])^(data_in[198]&H_in[2246])^(data_in[199]&H_in[2247])^(data_in[200]&H_in[2248])^(data_in[201]&H_in[2249])^(data_in[202]&H_in[2250])^(data_in[203]&H_in[2251])^(data_in[204]&H_in[2252])^(data_in[205]&H_in[2253])^(data_in[206]&H_in[2254])^(data_in[207]&H_in[2255])^(data_in[208]&H_in[2256])^(data_in[209]&H_in[2257])^(data_in[210]&H_in[2258])^(data_in[211]&H_in[2259])^(data_in[212]&H_in[2260])^(data_in[213]&H_in[2261])^(data_in[214]&H_in[2262])^(data_in[215]&H_in[2263])^(data_in[216]&H_in[2264])^(data_in[217]&H_in[2265])^(data_in[218]&H_in[2266])^(data_in[219]&H_in[2267])^(data_in[220]&H_in[2268])^(data_in[221]&H_in[2269])^(data_in[222]&H_in[2270])^(data_in[223]&H_in[2271])^(data_in[224]&H_in[2272])^(data_in[225]&H_in[2273])^(data_in[226]&H_in[2274])^(data_in[227]&H_in[2275])^(data_in[228]&H_in[2276])^(data_in[229]&H_in[2277])^(data_in[230]&H_in[2278])^(data_in[231]&H_in[2279])^(data_in[232]&H_in[2280])^(data_in[233]&H_in[2281])^(data_in[234]&H_in[2282])^(data_in[235]&H_in[2283])^(data_in[236]&H_in[2284])^(data_in[237]&H_in[2285])^(data_in[238]&H_in[2286])^(data_in[239]&H_in[2287])^(data_in[240]&H_in[2288])^(data_in[241]&H_in[2289])^(data_in[242]&H_in[2290])^(data_in[243]&H_in[2291])^(data_in[244]&H_in[2292])^(data_in[245]&H_in[2293])^(data_in[246]&H_in[2294])^(data_in[247]&H_in[2295])^(data_in[248]&H_in[2296])^(data_in[249]&H_in[2297])^(data_in[250]&H_in[2298])^(data_in[251]&H_in[2299])^(data_in[252]&H_in[2300])^(data_in[253]&H_in[2301])^(data_in[254]&H_in[2302])^(data_in[255]&H_in[2303]);
         data_out[9]<=(data_in[0]&H_in[2304])^(data_in[1]&H_in[2305])^(data_in[2]&H_in[2306])^(data_in[3]&H_in[2307])^(data_in[4]&H_in[2308])^(data_in[5]&H_in[2309])^(data_in[6]&H_in[2310])^(data_in[7]&H_in[2311])^(data_in[8]&H_in[2312])^(data_in[9]&H_in[2313])^(data_in[10]&H_in[2314])^(data_in[11]&H_in[2315])^(data_in[12]&H_in[2316])^(data_in[13]&H_in[2317])^(data_in[14]&H_in[2318])^(data_in[15]&H_in[2319])^(data_in[16]&H_in[2320])^(data_in[17]&H_in[2321])^(data_in[18]&H_in[2322])^(data_in[19]&H_in[2323])^(data_in[20]&H_in[2324])^(data_in[21]&H_in[2325])^(data_in[22]&H_in[2326])^(data_in[23]&H_in[2327])^(data_in[24]&H_in[2328])^(data_in[25]&H_in[2329])^(data_in[26]&H_in[2330])^(data_in[27]&H_in[2331])^(data_in[28]&H_in[2332])^(data_in[29]&H_in[2333])^(data_in[30]&H_in[2334])^(data_in[31]&H_in[2335])^(data_in[32]&H_in[2336])^(data_in[33]&H_in[2337])^(data_in[34]&H_in[2338])^(data_in[35]&H_in[2339])^(data_in[36]&H_in[2340])^(data_in[37]&H_in[2341])^(data_in[38]&H_in[2342])^(data_in[39]&H_in[2343])^(data_in[40]&H_in[2344])^(data_in[41]&H_in[2345])^(data_in[42]&H_in[2346])^(data_in[43]&H_in[2347])^(data_in[44]&H_in[2348])^(data_in[45]&H_in[2349])^(data_in[46]&H_in[2350])^(data_in[47]&H_in[2351])^(data_in[48]&H_in[2352])^(data_in[49]&H_in[2353])^(data_in[50]&H_in[2354])^(data_in[51]&H_in[2355])^(data_in[52]&H_in[2356])^(data_in[53]&H_in[2357])^(data_in[54]&H_in[2358])^(data_in[55]&H_in[2359])^(data_in[56]&H_in[2360])^(data_in[57]&H_in[2361])^(data_in[58]&H_in[2362])^(data_in[59]&H_in[2363])^(data_in[60]&H_in[2364])^(data_in[61]&H_in[2365])^(data_in[62]&H_in[2366])^(data_in[63]&H_in[2367])^(data_in[64]&H_in[2368])^(data_in[65]&H_in[2369])^(data_in[66]&H_in[2370])^(data_in[67]&H_in[2371])^(data_in[68]&H_in[2372])^(data_in[69]&H_in[2373])^(data_in[70]&H_in[2374])^(data_in[71]&H_in[2375])^(data_in[72]&H_in[2376])^(data_in[73]&H_in[2377])^(data_in[74]&H_in[2378])^(data_in[75]&H_in[2379])^(data_in[76]&H_in[2380])^(data_in[77]&H_in[2381])^(data_in[78]&H_in[2382])^(data_in[79]&H_in[2383])^(data_in[80]&H_in[2384])^(data_in[81]&H_in[2385])^(data_in[82]&H_in[2386])^(data_in[83]&H_in[2387])^(data_in[84]&H_in[2388])^(data_in[85]&H_in[2389])^(data_in[86]&H_in[2390])^(data_in[87]&H_in[2391])^(data_in[88]&H_in[2392])^(data_in[89]&H_in[2393])^(data_in[90]&H_in[2394])^(data_in[91]&H_in[2395])^(data_in[92]&H_in[2396])^(data_in[93]&H_in[2397])^(data_in[94]&H_in[2398])^(data_in[95]&H_in[2399])^(data_in[96]&H_in[2400])^(data_in[97]&H_in[2401])^(data_in[98]&H_in[2402])^(data_in[99]&H_in[2403])^(data_in[100]&H_in[2404])^(data_in[101]&H_in[2405])^(data_in[102]&H_in[2406])^(data_in[103]&H_in[2407])^(data_in[104]&H_in[2408])^(data_in[105]&H_in[2409])^(data_in[106]&H_in[2410])^(data_in[107]&H_in[2411])^(data_in[108]&H_in[2412])^(data_in[109]&H_in[2413])^(data_in[110]&H_in[2414])^(data_in[111]&H_in[2415])^(data_in[112]&H_in[2416])^(data_in[113]&H_in[2417])^(data_in[114]&H_in[2418])^(data_in[115]&H_in[2419])^(data_in[116]&H_in[2420])^(data_in[117]&H_in[2421])^(data_in[118]&H_in[2422])^(data_in[119]&H_in[2423])^(data_in[120]&H_in[2424])^(data_in[121]&H_in[2425])^(data_in[122]&H_in[2426])^(data_in[123]&H_in[2427])^(data_in[124]&H_in[2428])^(data_in[125]&H_in[2429])^(data_in[126]&H_in[2430])^(data_in[127]&H_in[2431])^(data_in[128]&H_in[2432])^(data_in[129]&H_in[2433])^(data_in[130]&H_in[2434])^(data_in[131]&H_in[2435])^(data_in[132]&H_in[2436])^(data_in[133]&H_in[2437])^(data_in[134]&H_in[2438])^(data_in[135]&H_in[2439])^(data_in[136]&H_in[2440])^(data_in[137]&H_in[2441])^(data_in[138]&H_in[2442])^(data_in[139]&H_in[2443])^(data_in[140]&H_in[2444])^(data_in[141]&H_in[2445])^(data_in[142]&H_in[2446])^(data_in[143]&H_in[2447])^(data_in[144]&H_in[2448])^(data_in[145]&H_in[2449])^(data_in[146]&H_in[2450])^(data_in[147]&H_in[2451])^(data_in[148]&H_in[2452])^(data_in[149]&H_in[2453])^(data_in[150]&H_in[2454])^(data_in[151]&H_in[2455])^(data_in[152]&H_in[2456])^(data_in[153]&H_in[2457])^(data_in[154]&H_in[2458])^(data_in[155]&H_in[2459])^(data_in[156]&H_in[2460])^(data_in[157]&H_in[2461])^(data_in[158]&H_in[2462])^(data_in[159]&H_in[2463])^(data_in[160]&H_in[2464])^(data_in[161]&H_in[2465])^(data_in[162]&H_in[2466])^(data_in[163]&H_in[2467])^(data_in[164]&H_in[2468])^(data_in[165]&H_in[2469])^(data_in[166]&H_in[2470])^(data_in[167]&H_in[2471])^(data_in[168]&H_in[2472])^(data_in[169]&H_in[2473])^(data_in[170]&H_in[2474])^(data_in[171]&H_in[2475])^(data_in[172]&H_in[2476])^(data_in[173]&H_in[2477])^(data_in[174]&H_in[2478])^(data_in[175]&H_in[2479])^(data_in[176]&H_in[2480])^(data_in[177]&H_in[2481])^(data_in[178]&H_in[2482])^(data_in[179]&H_in[2483])^(data_in[180]&H_in[2484])^(data_in[181]&H_in[2485])^(data_in[182]&H_in[2486])^(data_in[183]&H_in[2487])^(data_in[184]&H_in[2488])^(data_in[185]&H_in[2489])^(data_in[186]&H_in[2490])^(data_in[187]&H_in[2491])^(data_in[188]&H_in[2492])^(data_in[189]&H_in[2493])^(data_in[190]&H_in[2494])^(data_in[191]&H_in[2495])^(data_in[192]&H_in[2496])^(data_in[193]&H_in[2497])^(data_in[194]&H_in[2498])^(data_in[195]&H_in[2499])^(data_in[196]&H_in[2500])^(data_in[197]&H_in[2501])^(data_in[198]&H_in[2502])^(data_in[199]&H_in[2503])^(data_in[200]&H_in[2504])^(data_in[201]&H_in[2505])^(data_in[202]&H_in[2506])^(data_in[203]&H_in[2507])^(data_in[204]&H_in[2508])^(data_in[205]&H_in[2509])^(data_in[206]&H_in[2510])^(data_in[207]&H_in[2511])^(data_in[208]&H_in[2512])^(data_in[209]&H_in[2513])^(data_in[210]&H_in[2514])^(data_in[211]&H_in[2515])^(data_in[212]&H_in[2516])^(data_in[213]&H_in[2517])^(data_in[214]&H_in[2518])^(data_in[215]&H_in[2519])^(data_in[216]&H_in[2520])^(data_in[217]&H_in[2521])^(data_in[218]&H_in[2522])^(data_in[219]&H_in[2523])^(data_in[220]&H_in[2524])^(data_in[221]&H_in[2525])^(data_in[222]&H_in[2526])^(data_in[223]&H_in[2527])^(data_in[224]&H_in[2528])^(data_in[225]&H_in[2529])^(data_in[226]&H_in[2530])^(data_in[227]&H_in[2531])^(data_in[228]&H_in[2532])^(data_in[229]&H_in[2533])^(data_in[230]&H_in[2534])^(data_in[231]&H_in[2535])^(data_in[232]&H_in[2536])^(data_in[233]&H_in[2537])^(data_in[234]&H_in[2538])^(data_in[235]&H_in[2539])^(data_in[236]&H_in[2540])^(data_in[237]&H_in[2541])^(data_in[238]&H_in[2542])^(data_in[239]&H_in[2543])^(data_in[240]&H_in[2544])^(data_in[241]&H_in[2545])^(data_in[242]&H_in[2546])^(data_in[243]&H_in[2547])^(data_in[244]&H_in[2548])^(data_in[245]&H_in[2549])^(data_in[246]&H_in[2550])^(data_in[247]&H_in[2551])^(data_in[248]&H_in[2552])^(data_in[249]&H_in[2553])^(data_in[250]&H_in[2554])^(data_in[251]&H_in[2555])^(data_in[252]&H_in[2556])^(data_in[253]&H_in[2557])^(data_in[254]&H_in[2558])^(data_in[255]&H_in[2559]);
         data_out[10]<=(data_in[0]&H_in[2560])^(data_in[1]&H_in[2561])^(data_in[2]&H_in[2562])^(data_in[3]&H_in[2563])^(data_in[4]&H_in[2564])^(data_in[5]&H_in[2565])^(data_in[6]&H_in[2566])^(data_in[7]&H_in[2567])^(data_in[8]&H_in[2568])^(data_in[9]&H_in[2569])^(data_in[10]&H_in[2570])^(data_in[11]&H_in[2571])^(data_in[12]&H_in[2572])^(data_in[13]&H_in[2573])^(data_in[14]&H_in[2574])^(data_in[15]&H_in[2575])^(data_in[16]&H_in[2576])^(data_in[17]&H_in[2577])^(data_in[18]&H_in[2578])^(data_in[19]&H_in[2579])^(data_in[20]&H_in[2580])^(data_in[21]&H_in[2581])^(data_in[22]&H_in[2582])^(data_in[23]&H_in[2583])^(data_in[24]&H_in[2584])^(data_in[25]&H_in[2585])^(data_in[26]&H_in[2586])^(data_in[27]&H_in[2587])^(data_in[28]&H_in[2588])^(data_in[29]&H_in[2589])^(data_in[30]&H_in[2590])^(data_in[31]&H_in[2591])^(data_in[32]&H_in[2592])^(data_in[33]&H_in[2593])^(data_in[34]&H_in[2594])^(data_in[35]&H_in[2595])^(data_in[36]&H_in[2596])^(data_in[37]&H_in[2597])^(data_in[38]&H_in[2598])^(data_in[39]&H_in[2599])^(data_in[40]&H_in[2600])^(data_in[41]&H_in[2601])^(data_in[42]&H_in[2602])^(data_in[43]&H_in[2603])^(data_in[44]&H_in[2604])^(data_in[45]&H_in[2605])^(data_in[46]&H_in[2606])^(data_in[47]&H_in[2607])^(data_in[48]&H_in[2608])^(data_in[49]&H_in[2609])^(data_in[50]&H_in[2610])^(data_in[51]&H_in[2611])^(data_in[52]&H_in[2612])^(data_in[53]&H_in[2613])^(data_in[54]&H_in[2614])^(data_in[55]&H_in[2615])^(data_in[56]&H_in[2616])^(data_in[57]&H_in[2617])^(data_in[58]&H_in[2618])^(data_in[59]&H_in[2619])^(data_in[60]&H_in[2620])^(data_in[61]&H_in[2621])^(data_in[62]&H_in[2622])^(data_in[63]&H_in[2623])^(data_in[64]&H_in[2624])^(data_in[65]&H_in[2625])^(data_in[66]&H_in[2626])^(data_in[67]&H_in[2627])^(data_in[68]&H_in[2628])^(data_in[69]&H_in[2629])^(data_in[70]&H_in[2630])^(data_in[71]&H_in[2631])^(data_in[72]&H_in[2632])^(data_in[73]&H_in[2633])^(data_in[74]&H_in[2634])^(data_in[75]&H_in[2635])^(data_in[76]&H_in[2636])^(data_in[77]&H_in[2637])^(data_in[78]&H_in[2638])^(data_in[79]&H_in[2639])^(data_in[80]&H_in[2640])^(data_in[81]&H_in[2641])^(data_in[82]&H_in[2642])^(data_in[83]&H_in[2643])^(data_in[84]&H_in[2644])^(data_in[85]&H_in[2645])^(data_in[86]&H_in[2646])^(data_in[87]&H_in[2647])^(data_in[88]&H_in[2648])^(data_in[89]&H_in[2649])^(data_in[90]&H_in[2650])^(data_in[91]&H_in[2651])^(data_in[92]&H_in[2652])^(data_in[93]&H_in[2653])^(data_in[94]&H_in[2654])^(data_in[95]&H_in[2655])^(data_in[96]&H_in[2656])^(data_in[97]&H_in[2657])^(data_in[98]&H_in[2658])^(data_in[99]&H_in[2659])^(data_in[100]&H_in[2660])^(data_in[101]&H_in[2661])^(data_in[102]&H_in[2662])^(data_in[103]&H_in[2663])^(data_in[104]&H_in[2664])^(data_in[105]&H_in[2665])^(data_in[106]&H_in[2666])^(data_in[107]&H_in[2667])^(data_in[108]&H_in[2668])^(data_in[109]&H_in[2669])^(data_in[110]&H_in[2670])^(data_in[111]&H_in[2671])^(data_in[112]&H_in[2672])^(data_in[113]&H_in[2673])^(data_in[114]&H_in[2674])^(data_in[115]&H_in[2675])^(data_in[116]&H_in[2676])^(data_in[117]&H_in[2677])^(data_in[118]&H_in[2678])^(data_in[119]&H_in[2679])^(data_in[120]&H_in[2680])^(data_in[121]&H_in[2681])^(data_in[122]&H_in[2682])^(data_in[123]&H_in[2683])^(data_in[124]&H_in[2684])^(data_in[125]&H_in[2685])^(data_in[126]&H_in[2686])^(data_in[127]&H_in[2687])^(data_in[128]&H_in[2688])^(data_in[129]&H_in[2689])^(data_in[130]&H_in[2690])^(data_in[131]&H_in[2691])^(data_in[132]&H_in[2692])^(data_in[133]&H_in[2693])^(data_in[134]&H_in[2694])^(data_in[135]&H_in[2695])^(data_in[136]&H_in[2696])^(data_in[137]&H_in[2697])^(data_in[138]&H_in[2698])^(data_in[139]&H_in[2699])^(data_in[140]&H_in[2700])^(data_in[141]&H_in[2701])^(data_in[142]&H_in[2702])^(data_in[143]&H_in[2703])^(data_in[144]&H_in[2704])^(data_in[145]&H_in[2705])^(data_in[146]&H_in[2706])^(data_in[147]&H_in[2707])^(data_in[148]&H_in[2708])^(data_in[149]&H_in[2709])^(data_in[150]&H_in[2710])^(data_in[151]&H_in[2711])^(data_in[152]&H_in[2712])^(data_in[153]&H_in[2713])^(data_in[154]&H_in[2714])^(data_in[155]&H_in[2715])^(data_in[156]&H_in[2716])^(data_in[157]&H_in[2717])^(data_in[158]&H_in[2718])^(data_in[159]&H_in[2719])^(data_in[160]&H_in[2720])^(data_in[161]&H_in[2721])^(data_in[162]&H_in[2722])^(data_in[163]&H_in[2723])^(data_in[164]&H_in[2724])^(data_in[165]&H_in[2725])^(data_in[166]&H_in[2726])^(data_in[167]&H_in[2727])^(data_in[168]&H_in[2728])^(data_in[169]&H_in[2729])^(data_in[170]&H_in[2730])^(data_in[171]&H_in[2731])^(data_in[172]&H_in[2732])^(data_in[173]&H_in[2733])^(data_in[174]&H_in[2734])^(data_in[175]&H_in[2735])^(data_in[176]&H_in[2736])^(data_in[177]&H_in[2737])^(data_in[178]&H_in[2738])^(data_in[179]&H_in[2739])^(data_in[180]&H_in[2740])^(data_in[181]&H_in[2741])^(data_in[182]&H_in[2742])^(data_in[183]&H_in[2743])^(data_in[184]&H_in[2744])^(data_in[185]&H_in[2745])^(data_in[186]&H_in[2746])^(data_in[187]&H_in[2747])^(data_in[188]&H_in[2748])^(data_in[189]&H_in[2749])^(data_in[190]&H_in[2750])^(data_in[191]&H_in[2751])^(data_in[192]&H_in[2752])^(data_in[193]&H_in[2753])^(data_in[194]&H_in[2754])^(data_in[195]&H_in[2755])^(data_in[196]&H_in[2756])^(data_in[197]&H_in[2757])^(data_in[198]&H_in[2758])^(data_in[199]&H_in[2759])^(data_in[200]&H_in[2760])^(data_in[201]&H_in[2761])^(data_in[202]&H_in[2762])^(data_in[203]&H_in[2763])^(data_in[204]&H_in[2764])^(data_in[205]&H_in[2765])^(data_in[206]&H_in[2766])^(data_in[207]&H_in[2767])^(data_in[208]&H_in[2768])^(data_in[209]&H_in[2769])^(data_in[210]&H_in[2770])^(data_in[211]&H_in[2771])^(data_in[212]&H_in[2772])^(data_in[213]&H_in[2773])^(data_in[214]&H_in[2774])^(data_in[215]&H_in[2775])^(data_in[216]&H_in[2776])^(data_in[217]&H_in[2777])^(data_in[218]&H_in[2778])^(data_in[219]&H_in[2779])^(data_in[220]&H_in[2780])^(data_in[221]&H_in[2781])^(data_in[222]&H_in[2782])^(data_in[223]&H_in[2783])^(data_in[224]&H_in[2784])^(data_in[225]&H_in[2785])^(data_in[226]&H_in[2786])^(data_in[227]&H_in[2787])^(data_in[228]&H_in[2788])^(data_in[229]&H_in[2789])^(data_in[230]&H_in[2790])^(data_in[231]&H_in[2791])^(data_in[232]&H_in[2792])^(data_in[233]&H_in[2793])^(data_in[234]&H_in[2794])^(data_in[235]&H_in[2795])^(data_in[236]&H_in[2796])^(data_in[237]&H_in[2797])^(data_in[238]&H_in[2798])^(data_in[239]&H_in[2799])^(data_in[240]&H_in[2800])^(data_in[241]&H_in[2801])^(data_in[242]&H_in[2802])^(data_in[243]&H_in[2803])^(data_in[244]&H_in[2804])^(data_in[245]&H_in[2805])^(data_in[246]&H_in[2806])^(data_in[247]&H_in[2807])^(data_in[248]&H_in[2808])^(data_in[249]&H_in[2809])^(data_in[250]&H_in[2810])^(data_in[251]&H_in[2811])^(data_in[252]&H_in[2812])^(data_in[253]&H_in[2813])^(data_in[254]&H_in[2814])^(data_in[255]&H_in[2815]);
         data_out[11]<=(data_in[0]&H_in[2816])^(data_in[1]&H_in[2817])^(data_in[2]&H_in[2818])^(data_in[3]&H_in[2819])^(data_in[4]&H_in[2820])^(data_in[5]&H_in[2821])^(data_in[6]&H_in[2822])^(data_in[7]&H_in[2823])^(data_in[8]&H_in[2824])^(data_in[9]&H_in[2825])^(data_in[10]&H_in[2826])^(data_in[11]&H_in[2827])^(data_in[12]&H_in[2828])^(data_in[13]&H_in[2829])^(data_in[14]&H_in[2830])^(data_in[15]&H_in[2831])^(data_in[16]&H_in[2832])^(data_in[17]&H_in[2833])^(data_in[18]&H_in[2834])^(data_in[19]&H_in[2835])^(data_in[20]&H_in[2836])^(data_in[21]&H_in[2837])^(data_in[22]&H_in[2838])^(data_in[23]&H_in[2839])^(data_in[24]&H_in[2840])^(data_in[25]&H_in[2841])^(data_in[26]&H_in[2842])^(data_in[27]&H_in[2843])^(data_in[28]&H_in[2844])^(data_in[29]&H_in[2845])^(data_in[30]&H_in[2846])^(data_in[31]&H_in[2847])^(data_in[32]&H_in[2848])^(data_in[33]&H_in[2849])^(data_in[34]&H_in[2850])^(data_in[35]&H_in[2851])^(data_in[36]&H_in[2852])^(data_in[37]&H_in[2853])^(data_in[38]&H_in[2854])^(data_in[39]&H_in[2855])^(data_in[40]&H_in[2856])^(data_in[41]&H_in[2857])^(data_in[42]&H_in[2858])^(data_in[43]&H_in[2859])^(data_in[44]&H_in[2860])^(data_in[45]&H_in[2861])^(data_in[46]&H_in[2862])^(data_in[47]&H_in[2863])^(data_in[48]&H_in[2864])^(data_in[49]&H_in[2865])^(data_in[50]&H_in[2866])^(data_in[51]&H_in[2867])^(data_in[52]&H_in[2868])^(data_in[53]&H_in[2869])^(data_in[54]&H_in[2870])^(data_in[55]&H_in[2871])^(data_in[56]&H_in[2872])^(data_in[57]&H_in[2873])^(data_in[58]&H_in[2874])^(data_in[59]&H_in[2875])^(data_in[60]&H_in[2876])^(data_in[61]&H_in[2877])^(data_in[62]&H_in[2878])^(data_in[63]&H_in[2879])^(data_in[64]&H_in[2880])^(data_in[65]&H_in[2881])^(data_in[66]&H_in[2882])^(data_in[67]&H_in[2883])^(data_in[68]&H_in[2884])^(data_in[69]&H_in[2885])^(data_in[70]&H_in[2886])^(data_in[71]&H_in[2887])^(data_in[72]&H_in[2888])^(data_in[73]&H_in[2889])^(data_in[74]&H_in[2890])^(data_in[75]&H_in[2891])^(data_in[76]&H_in[2892])^(data_in[77]&H_in[2893])^(data_in[78]&H_in[2894])^(data_in[79]&H_in[2895])^(data_in[80]&H_in[2896])^(data_in[81]&H_in[2897])^(data_in[82]&H_in[2898])^(data_in[83]&H_in[2899])^(data_in[84]&H_in[2900])^(data_in[85]&H_in[2901])^(data_in[86]&H_in[2902])^(data_in[87]&H_in[2903])^(data_in[88]&H_in[2904])^(data_in[89]&H_in[2905])^(data_in[90]&H_in[2906])^(data_in[91]&H_in[2907])^(data_in[92]&H_in[2908])^(data_in[93]&H_in[2909])^(data_in[94]&H_in[2910])^(data_in[95]&H_in[2911])^(data_in[96]&H_in[2912])^(data_in[97]&H_in[2913])^(data_in[98]&H_in[2914])^(data_in[99]&H_in[2915])^(data_in[100]&H_in[2916])^(data_in[101]&H_in[2917])^(data_in[102]&H_in[2918])^(data_in[103]&H_in[2919])^(data_in[104]&H_in[2920])^(data_in[105]&H_in[2921])^(data_in[106]&H_in[2922])^(data_in[107]&H_in[2923])^(data_in[108]&H_in[2924])^(data_in[109]&H_in[2925])^(data_in[110]&H_in[2926])^(data_in[111]&H_in[2927])^(data_in[112]&H_in[2928])^(data_in[113]&H_in[2929])^(data_in[114]&H_in[2930])^(data_in[115]&H_in[2931])^(data_in[116]&H_in[2932])^(data_in[117]&H_in[2933])^(data_in[118]&H_in[2934])^(data_in[119]&H_in[2935])^(data_in[120]&H_in[2936])^(data_in[121]&H_in[2937])^(data_in[122]&H_in[2938])^(data_in[123]&H_in[2939])^(data_in[124]&H_in[2940])^(data_in[125]&H_in[2941])^(data_in[126]&H_in[2942])^(data_in[127]&H_in[2943])^(data_in[128]&H_in[2944])^(data_in[129]&H_in[2945])^(data_in[130]&H_in[2946])^(data_in[131]&H_in[2947])^(data_in[132]&H_in[2948])^(data_in[133]&H_in[2949])^(data_in[134]&H_in[2950])^(data_in[135]&H_in[2951])^(data_in[136]&H_in[2952])^(data_in[137]&H_in[2953])^(data_in[138]&H_in[2954])^(data_in[139]&H_in[2955])^(data_in[140]&H_in[2956])^(data_in[141]&H_in[2957])^(data_in[142]&H_in[2958])^(data_in[143]&H_in[2959])^(data_in[144]&H_in[2960])^(data_in[145]&H_in[2961])^(data_in[146]&H_in[2962])^(data_in[147]&H_in[2963])^(data_in[148]&H_in[2964])^(data_in[149]&H_in[2965])^(data_in[150]&H_in[2966])^(data_in[151]&H_in[2967])^(data_in[152]&H_in[2968])^(data_in[153]&H_in[2969])^(data_in[154]&H_in[2970])^(data_in[155]&H_in[2971])^(data_in[156]&H_in[2972])^(data_in[157]&H_in[2973])^(data_in[158]&H_in[2974])^(data_in[159]&H_in[2975])^(data_in[160]&H_in[2976])^(data_in[161]&H_in[2977])^(data_in[162]&H_in[2978])^(data_in[163]&H_in[2979])^(data_in[164]&H_in[2980])^(data_in[165]&H_in[2981])^(data_in[166]&H_in[2982])^(data_in[167]&H_in[2983])^(data_in[168]&H_in[2984])^(data_in[169]&H_in[2985])^(data_in[170]&H_in[2986])^(data_in[171]&H_in[2987])^(data_in[172]&H_in[2988])^(data_in[173]&H_in[2989])^(data_in[174]&H_in[2990])^(data_in[175]&H_in[2991])^(data_in[176]&H_in[2992])^(data_in[177]&H_in[2993])^(data_in[178]&H_in[2994])^(data_in[179]&H_in[2995])^(data_in[180]&H_in[2996])^(data_in[181]&H_in[2997])^(data_in[182]&H_in[2998])^(data_in[183]&H_in[2999])^(data_in[184]&H_in[3000])^(data_in[185]&H_in[3001])^(data_in[186]&H_in[3002])^(data_in[187]&H_in[3003])^(data_in[188]&H_in[3004])^(data_in[189]&H_in[3005])^(data_in[190]&H_in[3006])^(data_in[191]&H_in[3007])^(data_in[192]&H_in[3008])^(data_in[193]&H_in[3009])^(data_in[194]&H_in[3010])^(data_in[195]&H_in[3011])^(data_in[196]&H_in[3012])^(data_in[197]&H_in[3013])^(data_in[198]&H_in[3014])^(data_in[199]&H_in[3015])^(data_in[200]&H_in[3016])^(data_in[201]&H_in[3017])^(data_in[202]&H_in[3018])^(data_in[203]&H_in[3019])^(data_in[204]&H_in[3020])^(data_in[205]&H_in[3021])^(data_in[206]&H_in[3022])^(data_in[207]&H_in[3023])^(data_in[208]&H_in[3024])^(data_in[209]&H_in[3025])^(data_in[210]&H_in[3026])^(data_in[211]&H_in[3027])^(data_in[212]&H_in[3028])^(data_in[213]&H_in[3029])^(data_in[214]&H_in[3030])^(data_in[215]&H_in[3031])^(data_in[216]&H_in[3032])^(data_in[217]&H_in[3033])^(data_in[218]&H_in[3034])^(data_in[219]&H_in[3035])^(data_in[220]&H_in[3036])^(data_in[221]&H_in[3037])^(data_in[222]&H_in[3038])^(data_in[223]&H_in[3039])^(data_in[224]&H_in[3040])^(data_in[225]&H_in[3041])^(data_in[226]&H_in[3042])^(data_in[227]&H_in[3043])^(data_in[228]&H_in[3044])^(data_in[229]&H_in[3045])^(data_in[230]&H_in[3046])^(data_in[231]&H_in[3047])^(data_in[232]&H_in[3048])^(data_in[233]&H_in[3049])^(data_in[234]&H_in[3050])^(data_in[235]&H_in[3051])^(data_in[236]&H_in[3052])^(data_in[237]&H_in[3053])^(data_in[238]&H_in[3054])^(data_in[239]&H_in[3055])^(data_in[240]&H_in[3056])^(data_in[241]&H_in[3057])^(data_in[242]&H_in[3058])^(data_in[243]&H_in[3059])^(data_in[244]&H_in[3060])^(data_in[245]&H_in[3061])^(data_in[246]&H_in[3062])^(data_in[247]&H_in[3063])^(data_in[248]&H_in[3064])^(data_in[249]&H_in[3065])^(data_in[250]&H_in[3066])^(data_in[251]&H_in[3067])^(data_in[252]&H_in[3068])^(data_in[253]&H_in[3069])^(data_in[254]&H_in[3070])^(data_in[255]&H_in[3071]);
         data_out[12]<=(data_in[0]&H_in[3072])^(data_in[1]&H_in[3073])^(data_in[2]&H_in[3074])^(data_in[3]&H_in[3075])^(data_in[4]&H_in[3076])^(data_in[5]&H_in[3077])^(data_in[6]&H_in[3078])^(data_in[7]&H_in[3079])^(data_in[8]&H_in[3080])^(data_in[9]&H_in[3081])^(data_in[10]&H_in[3082])^(data_in[11]&H_in[3083])^(data_in[12]&H_in[3084])^(data_in[13]&H_in[3085])^(data_in[14]&H_in[3086])^(data_in[15]&H_in[3087])^(data_in[16]&H_in[3088])^(data_in[17]&H_in[3089])^(data_in[18]&H_in[3090])^(data_in[19]&H_in[3091])^(data_in[20]&H_in[3092])^(data_in[21]&H_in[3093])^(data_in[22]&H_in[3094])^(data_in[23]&H_in[3095])^(data_in[24]&H_in[3096])^(data_in[25]&H_in[3097])^(data_in[26]&H_in[3098])^(data_in[27]&H_in[3099])^(data_in[28]&H_in[3100])^(data_in[29]&H_in[3101])^(data_in[30]&H_in[3102])^(data_in[31]&H_in[3103])^(data_in[32]&H_in[3104])^(data_in[33]&H_in[3105])^(data_in[34]&H_in[3106])^(data_in[35]&H_in[3107])^(data_in[36]&H_in[3108])^(data_in[37]&H_in[3109])^(data_in[38]&H_in[3110])^(data_in[39]&H_in[3111])^(data_in[40]&H_in[3112])^(data_in[41]&H_in[3113])^(data_in[42]&H_in[3114])^(data_in[43]&H_in[3115])^(data_in[44]&H_in[3116])^(data_in[45]&H_in[3117])^(data_in[46]&H_in[3118])^(data_in[47]&H_in[3119])^(data_in[48]&H_in[3120])^(data_in[49]&H_in[3121])^(data_in[50]&H_in[3122])^(data_in[51]&H_in[3123])^(data_in[52]&H_in[3124])^(data_in[53]&H_in[3125])^(data_in[54]&H_in[3126])^(data_in[55]&H_in[3127])^(data_in[56]&H_in[3128])^(data_in[57]&H_in[3129])^(data_in[58]&H_in[3130])^(data_in[59]&H_in[3131])^(data_in[60]&H_in[3132])^(data_in[61]&H_in[3133])^(data_in[62]&H_in[3134])^(data_in[63]&H_in[3135])^(data_in[64]&H_in[3136])^(data_in[65]&H_in[3137])^(data_in[66]&H_in[3138])^(data_in[67]&H_in[3139])^(data_in[68]&H_in[3140])^(data_in[69]&H_in[3141])^(data_in[70]&H_in[3142])^(data_in[71]&H_in[3143])^(data_in[72]&H_in[3144])^(data_in[73]&H_in[3145])^(data_in[74]&H_in[3146])^(data_in[75]&H_in[3147])^(data_in[76]&H_in[3148])^(data_in[77]&H_in[3149])^(data_in[78]&H_in[3150])^(data_in[79]&H_in[3151])^(data_in[80]&H_in[3152])^(data_in[81]&H_in[3153])^(data_in[82]&H_in[3154])^(data_in[83]&H_in[3155])^(data_in[84]&H_in[3156])^(data_in[85]&H_in[3157])^(data_in[86]&H_in[3158])^(data_in[87]&H_in[3159])^(data_in[88]&H_in[3160])^(data_in[89]&H_in[3161])^(data_in[90]&H_in[3162])^(data_in[91]&H_in[3163])^(data_in[92]&H_in[3164])^(data_in[93]&H_in[3165])^(data_in[94]&H_in[3166])^(data_in[95]&H_in[3167])^(data_in[96]&H_in[3168])^(data_in[97]&H_in[3169])^(data_in[98]&H_in[3170])^(data_in[99]&H_in[3171])^(data_in[100]&H_in[3172])^(data_in[101]&H_in[3173])^(data_in[102]&H_in[3174])^(data_in[103]&H_in[3175])^(data_in[104]&H_in[3176])^(data_in[105]&H_in[3177])^(data_in[106]&H_in[3178])^(data_in[107]&H_in[3179])^(data_in[108]&H_in[3180])^(data_in[109]&H_in[3181])^(data_in[110]&H_in[3182])^(data_in[111]&H_in[3183])^(data_in[112]&H_in[3184])^(data_in[113]&H_in[3185])^(data_in[114]&H_in[3186])^(data_in[115]&H_in[3187])^(data_in[116]&H_in[3188])^(data_in[117]&H_in[3189])^(data_in[118]&H_in[3190])^(data_in[119]&H_in[3191])^(data_in[120]&H_in[3192])^(data_in[121]&H_in[3193])^(data_in[122]&H_in[3194])^(data_in[123]&H_in[3195])^(data_in[124]&H_in[3196])^(data_in[125]&H_in[3197])^(data_in[126]&H_in[3198])^(data_in[127]&H_in[3199])^(data_in[128]&H_in[3200])^(data_in[129]&H_in[3201])^(data_in[130]&H_in[3202])^(data_in[131]&H_in[3203])^(data_in[132]&H_in[3204])^(data_in[133]&H_in[3205])^(data_in[134]&H_in[3206])^(data_in[135]&H_in[3207])^(data_in[136]&H_in[3208])^(data_in[137]&H_in[3209])^(data_in[138]&H_in[3210])^(data_in[139]&H_in[3211])^(data_in[140]&H_in[3212])^(data_in[141]&H_in[3213])^(data_in[142]&H_in[3214])^(data_in[143]&H_in[3215])^(data_in[144]&H_in[3216])^(data_in[145]&H_in[3217])^(data_in[146]&H_in[3218])^(data_in[147]&H_in[3219])^(data_in[148]&H_in[3220])^(data_in[149]&H_in[3221])^(data_in[150]&H_in[3222])^(data_in[151]&H_in[3223])^(data_in[152]&H_in[3224])^(data_in[153]&H_in[3225])^(data_in[154]&H_in[3226])^(data_in[155]&H_in[3227])^(data_in[156]&H_in[3228])^(data_in[157]&H_in[3229])^(data_in[158]&H_in[3230])^(data_in[159]&H_in[3231])^(data_in[160]&H_in[3232])^(data_in[161]&H_in[3233])^(data_in[162]&H_in[3234])^(data_in[163]&H_in[3235])^(data_in[164]&H_in[3236])^(data_in[165]&H_in[3237])^(data_in[166]&H_in[3238])^(data_in[167]&H_in[3239])^(data_in[168]&H_in[3240])^(data_in[169]&H_in[3241])^(data_in[170]&H_in[3242])^(data_in[171]&H_in[3243])^(data_in[172]&H_in[3244])^(data_in[173]&H_in[3245])^(data_in[174]&H_in[3246])^(data_in[175]&H_in[3247])^(data_in[176]&H_in[3248])^(data_in[177]&H_in[3249])^(data_in[178]&H_in[3250])^(data_in[179]&H_in[3251])^(data_in[180]&H_in[3252])^(data_in[181]&H_in[3253])^(data_in[182]&H_in[3254])^(data_in[183]&H_in[3255])^(data_in[184]&H_in[3256])^(data_in[185]&H_in[3257])^(data_in[186]&H_in[3258])^(data_in[187]&H_in[3259])^(data_in[188]&H_in[3260])^(data_in[189]&H_in[3261])^(data_in[190]&H_in[3262])^(data_in[191]&H_in[3263])^(data_in[192]&H_in[3264])^(data_in[193]&H_in[3265])^(data_in[194]&H_in[3266])^(data_in[195]&H_in[3267])^(data_in[196]&H_in[3268])^(data_in[197]&H_in[3269])^(data_in[198]&H_in[3270])^(data_in[199]&H_in[3271])^(data_in[200]&H_in[3272])^(data_in[201]&H_in[3273])^(data_in[202]&H_in[3274])^(data_in[203]&H_in[3275])^(data_in[204]&H_in[3276])^(data_in[205]&H_in[3277])^(data_in[206]&H_in[3278])^(data_in[207]&H_in[3279])^(data_in[208]&H_in[3280])^(data_in[209]&H_in[3281])^(data_in[210]&H_in[3282])^(data_in[211]&H_in[3283])^(data_in[212]&H_in[3284])^(data_in[213]&H_in[3285])^(data_in[214]&H_in[3286])^(data_in[215]&H_in[3287])^(data_in[216]&H_in[3288])^(data_in[217]&H_in[3289])^(data_in[218]&H_in[3290])^(data_in[219]&H_in[3291])^(data_in[220]&H_in[3292])^(data_in[221]&H_in[3293])^(data_in[222]&H_in[3294])^(data_in[223]&H_in[3295])^(data_in[224]&H_in[3296])^(data_in[225]&H_in[3297])^(data_in[226]&H_in[3298])^(data_in[227]&H_in[3299])^(data_in[228]&H_in[3300])^(data_in[229]&H_in[3301])^(data_in[230]&H_in[3302])^(data_in[231]&H_in[3303])^(data_in[232]&H_in[3304])^(data_in[233]&H_in[3305])^(data_in[234]&H_in[3306])^(data_in[235]&H_in[3307])^(data_in[236]&H_in[3308])^(data_in[237]&H_in[3309])^(data_in[238]&H_in[3310])^(data_in[239]&H_in[3311])^(data_in[240]&H_in[3312])^(data_in[241]&H_in[3313])^(data_in[242]&H_in[3314])^(data_in[243]&H_in[3315])^(data_in[244]&H_in[3316])^(data_in[245]&H_in[3317])^(data_in[246]&H_in[3318])^(data_in[247]&H_in[3319])^(data_in[248]&H_in[3320])^(data_in[249]&H_in[3321])^(data_in[250]&H_in[3322])^(data_in[251]&H_in[3323])^(data_in[252]&H_in[3324])^(data_in[253]&H_in[3325])^(data_in[254]&H_in[3326])^(data_in[255]&H_in[3327]);
         data_out[13]<=(data_in[0]&H_in[3328])^(data_in[1]&H_in[3329])^(data_in[2]&H_in[3330])^(data_in[3]&H_in[3331])^(data_in[4]&H_in[3332])^(data_in[5]&H_in[3333])^(data_in[6]&H_in[3334])^(data_in[7]&H_in[3335])^(data_in[8]&H_in[3336])^(data_in[9]&H_in[3337])^(data_in[10]&H_in[3338])^(data_in[11]&H_in[3339])^(data_in[12]&H_in[3340])^(data_in[13]&H_in[3341])^(data_in[14]&H_in[3342])^(data_in[15]&H_in[3343])^(data_in[16]&H_in[3344])^(data_in[17]&H_in[3345])^(data_in[18]&H_in[3346])^(data_in[19]&H_in[3347])^(data_in[20]&H_in[3348])^(data_in[21]&H_in[3349])^(data_in[22]&H_in[3350])^(data_in[23]&H_in[3351])^(data_in[24]&H_in[3352])^(data_in[25]&H_in[3353])^(data_in[26]&H_in[3354])^(data_in[27]&H_in[3355])^(data_in[28]&H_in[3356])^(data_in[29]&H_in[3357])^(data_in[30]&H_in[3358])^(data_in[31]&H_in[3359])^(data_in[32]&H_in[3360])^(data_in[33]&H_in[3361])^(data_in[34]&H_in[3362])^(data_in[35]&H_in[3363])^(data_in[36]&H_in[3364])^(data_in[37]&H_in[3365])^(data_in[38]&H_in[3366])^(data_in[39]&H_in[3367])^(data_in[40]&H_in[3368])^(data_in[41]&H_in[3369])^(data_in[42]&H_in[3370])^(data_in[43]&H_in[3371])^(data_in[44]&H_in[3372])^(data_in[45]&H_in[3373])^(data_in[46]&H_in[3374])^(data_in[47]&H_in[3375])^(data_in[48]&H_in[3376])^(data_in[49]&H_in[3377])^(data_in[50]&H_in[3378])^(data_in[51]&H_in[3379])^(data_in[52]&H_in[3380])^(data_in[53]&H_in[3381])^(data_in[54]&H_in[3382])^(data_in[55]&H_in[3383])^(data_in[56]&H_in[3384])^(data_in[57]&H_in[3385])^(data_in[58]&H_in[3386])^(data_in[59]&H_in[3387])^(data_in[60]&H_in[3388])^(data_in[61]&H_in[3389])^(data_in[62]&H_in[3390])^(data_in[63]&H_in[3391])^(data_in[64]&H_in[3392])^(data_in[65]&H_in[3393])^(data_in[66]&H_in[3394])^(data_in[67]&H_in[3395])^(data_in[68]&H_in[3396])^(data_in[69]&H_in[3397])^(data_in[70]&H_in[3398])^(data_in[71]&H_in[3399])^(data_in[72]&H_in[3400])^(data_in[73]&H_in[3401])^(data_in[74]&H_in[3402])^(data_in[75]&H_in[3403])^(data_in[76]&H_in[3404])^(data_in[77]&H_in[3405])^(data_in[78]&H_in[3406])^(data_in[79]&H_in[3407])^(data_in[80]&H_in[3408])^(data_in[81]&H_in[3409])^(data_in[82]&H_in[3410])^(data_in[83]&H_in[3411])^(data_in[84]&H_in[3412])^(data_in[85]&H_in[3413])^(data_in[86]&H_in[3414])^(data_in[87]&H_in[3415])^(data_in[88]&H_in[3416])^(data_in[89]&H_in[3417])^(data_in[90]&H_in[3418])^(data_in[91]&H_in[3419])^(data_in[92]&H_in[3420])^(data_in[93]&H_in[3421])^(data_in[94]&H_in[3422])^(data_in[95]&H_in[3423])^(data_in[96]&H_in[3424])^(data_in[97]&H_in[3425])^(data_in[98]&H_in[3426])^(data_in[99]&H_in[3427])^(data_in[100]&H_in[3428])^(data_in[101]&H_in[3429])^(data_in[102]&H_in[3430])^(data_in[103]&H_in[3431])^(data_in[104]&H_in[3432])^(data_in[105]&H_in[3433])^(data_in[106]&H_in[3434])^(data_in[107]&H_in[3435])^(data_in[108]&H_in[3436])^(data_in[109]&H_in[3437])^(data_in[110]&H_in[3438])^(data_in[111]&H_in[3439])^(data_in[112]&H_in[3440])^(data_in[113]&H_in[3441])^(data_in[114]&H_in[3442])^(data_in[115]&H_in[3443])^(data_in[116]&H_in[3444])^(data_in[117]&H_in[3445])^(data_in[118]&H_in[3446])^(data_in[119]&H_in[3447])^(data_in[120]&H_in[3448])^(data_in[121]&H_in[3449])^(data_in[122]&H_in[3450])^(data_in[123]&H_in[3451])^(data_in[124]&H_in[3452])^(data_in[125]&H_in[3453])^(data_in[126]&H_in[3454])^(data_in[127]&H_in[3455])^(data_in[128]&H_in[3456])^(data_in[129]&H_in[3457])^(data_in[130]&H_in[3458])^(data_in[131]&H_in[3459])^(data_in[132]&H_in[3460])^(data_in[133]&H_in[3461])^(data_in[134]&H_in[3462])^(data_in[135]&H_in[3463])^(data_in[136]&H_in[3464])^(data_in[137]&H_in[3465])^(data_in[138]&H_in[3466])^(data_in[139]&H_in[3467])^(data_in[140]&H_in[3468])^(data_in[141]&H_in[3469])^(data_in[142]&H_in[3470])^(data_in[143]&H_in[3471])^(data_in[144]&H_in[3472])^(data_in[145]&H_in[3473])^(data_in[146]&H_in[3474])^(data_in[147]&H_in[3475])^(data_in[148]&H_in[3476])^(data_in[149]&H_in[3477])^(data_in[150]&H_in[3478])^(data_in[151]&H_in[3479])^(data_in[152]&H_in[3480])^(data_in[153]&H_in[3481])^(data_in[154]&H_in[3482])^(data_in[155]&H_in[3483])^(data_in[156]&H_in[3484])^(data_in[157]&H_in[3485])^(data_in[158]&H_in[3486])^(data_in[159]&H_in[3487])^(data_in[160]&H_in[3488])^(data_in[161]&H_in[3489])^(data_in[162]&H_in[3490])^(data_in[163]&H_in[3491])^(data_in[164]&H_in[3492])^(data_in[165]&H_in[3493])^(data_in[166]&H_in[3494])^(data_in[167]&H_in[3495])^(data_in[168]&H_in[3496])^(data_in[169]&H_in[3497])^(data_in[170]&H_in[3498])^(data_in[171]&H_in[3499])^(data_in[172]&H_in[3500])^(data_in[173]&H_in[3501])^(data_in[174]&H_in[3502])^(data_in[175]&H_in[3503])^(data_in[176]&H_in[3504])^(data_in[177]&H_in[3505])^(data_in[178]&H_in[3506])^(data_in[179]&H_in[3507])^(data_in[180]&H_in[3508])^(data_in[181]&H_in[3509])^(data_in[182]&H_in[3510])^(data_in[183]&H_in[3511])^(data_in[184]&H_in[3512])^(data_in[185]&H_in[3513])^(data_in[186]&H_in[3514])^(data_in[187]&H_in[3515])^(data_in[188]&H_in[3516])^(data_in[189]&H_in[3517])^(data_in[190]&H_in[3518])^(data_in[191]&H_in[3519])^(data_in[192]&H_in[3520])^(data_in[193]&H_in[3521])^(data_in[194]&H_in[3522])^(data_in[195]&H_in[3523])^(data_in[196]&H_in[3524])^(data_in[197]&H_in[3525])^(data_in[198]&H_in[3526])^(data_in[199]&H_in[3527])^(data_in[200]&H_in[3528])^(data_in[201]&H_in[3529])^(data_in[202]&H_in[3530])^(data_in[203]&H_in[3531])^(data_in[204]&H_in[3532])^(data_in[205]&H_in[3533])^(data_in[206]&H_in[3534])^(data_in[207]&H_in[3535])^(data_in[208]&H_in[3536])^(data_in[209]&H_in[3537])^(data_in[210]&H_in[3538])^(data_in[211]&H_in[3539])^(data_in[212]&H_in[3540])^(data_in[213]&H_in[3541])^(data_in[214]&H_in[3542])^(data_in[215]&H_in[3543])^(data_in[216]&H_in[3544])^(data_in[217]&H_in[3545])^(data_in[218]&H_in[3546])^(data_in[219]&H_in[3547])^(data_in[220]&H_in[3548])^(data_in[221]&H_in[3549])^(data_in[222]&H_in[3550])^(data_in[223]&H_in[3551])^(data_in[224]&H_in[3552])^(data_in[225]&H_in[3553])^(data_in[226]&H_in[3554])^(data_in[227]&H_in[3555])^(data_in[228]&H_in[3556])^(data_in[229]&H_in[3557])^(data_in[230]&H_in[3558])^(data_in[231]&H_in[3559])^(data_in[232]&H_in[3560])^(data_in[233]&H_in[3561])^(data_in[234]&H_in[3562])^(data_in[235]&H_in[3563])^(data_in[236]&H_in[3564])^(data_in[237]&H_in[3565])^(data_in[238]&H_in[3566])^(data_in[239]&H_in[3567])^(data_in[240]&H_in[3568])^(data_in[241]&H_in[3569])^(data_in[242]&H_in[3570])^(data_in[243]&H_in[3571])^(data_in[244]&H_in[3572])^(data_in[245]&H_in[3573])^(data_in[246]&H_in[3574])^(data_in[247]&H_in[3575])^(data_in[248]&H_in[3576])^(data_in[249]&H_in[3577])^(data_in[250]&H_in[3578])^(data_in[251]&H_in[3579])^(data_in[252]&H_in[3580])^(data_in[253]&H_in[3581])^(data_in[254]&H_in[3582])^(data_in[255]&H_in[3583]);
         data_out[14]<=(data_in[0]&H_in[3584])^(data_in[1]&H_in[3585])^(data_in[2]&H_in[3586])^(data_in[3]&H_in[3587])^(data_in[4]&H_in[3588])^(data_in[5]&H_in[3589])^(data_in[6]&H_in[3590])^(data_in[7]&H_in[3591])^(data_in[8]&H_in[3592])^(data_in[9]&H_in[3593])^(data_in[10]&H_in[3594])^(data_in[11]&H_in[3595])^(data_in[12]&H_in[3596])^(data_in[13]&H_in[3597])^(data_in[14]&H_in[3598])^(data_in[15]&H_in[3599])^(data_in[16]&H_in[3600])^(data_in[17]&H_in[3601])^(data_in[18]&H_in[3602])^(data_in[19]&H_in[3603])^(data_in[20]&H_in[3604])^(data_in[21]&H_in[3605])^(data_in[22]&H_in[3606])^(data_in[23]&H_in[3607])^(data_in[24]&H_in[3608])^(data_in[25]&H_in[3609])^(data_in[26]&H_in[3610])^(data_in[27]&H_in[3611])^(data_in[28]&H_in[3612])^(data_in[29]&H_in[3613])^(data_in[30]&H_in[3614])^(data_in[31]&H_in[3615])^(data_in[32]&H_in[3616])^(data_in[33]&H_in[3617])^(data_in[34]&H_in[3618])^(data_in[35]&H_in[3619])^(data_in[36]&H_in[3620])^(data_in[37]&H_in[3621])^(data_in[38]&H_in[3622])^(data_in[39]&H_in[3623])^(data_in[40]&H_in[3624])^(data_in[41]&H_in[3625])^(data_in[42]&H_in[3626])^(data_in[43]&H_in[3627])^(data_in[44]&H_in[3628])^(data_in[45]&H_in[3629])^(data_in[46]&H_in[3630])^(data_in[47]&H_in[3631])^(data_in[48]&H_in[3632])^(data_in[49]&H_in[3633])^(data_in[50]&H_in[3634])^(data_in[51]&H_in[3635])^(data_in[52]&H_in[3636])^(data_in[53]&H_in[3637])^(data_in[54]&H_in[3638])^(data_in[55]&H_in[3639])^(data_in[56]&H_in[3640])^(data_in[57]&H_in[3641])^(data_in[58]&H_in[3642])^(data_in[59]&H_in[3643])^(data_in[60]&H_in[3644])^(data_in[61]&H_in[3645])^(data_in[62]&H_in[3646])^(data_in[63]&H_in[3647])^(data_in[64]&H_in[3648])^(data_in[65]&H_in[3649])^(data_in[66]&H_in[3650])^(data_in[67]&H_in[3651])^(data_in[68]&H_in[3652])^(data_in[69]&H_in[3653])^(data_in[70]&H_in[3654])^(data_in[71]&H_in[3655])^(data_in[72]&H_in[3656])^(data_in[73]&H_in[3657])^(data_in[74]&H_in[3658])^(data_in[75]&H_in[3659])^(data_in[76]&H_in[3660])^(data_in[77]&H_in[3661])^(data_in[78]&H_in[3662])^(data_in[79]&H_in[3663])^(data_in[80]&H_in[3664])^(data_in[81]&H_in[3665])^(data_in[82]&H_in[3666])^(data_in[83]&H_in[3667])^(data_in[84]&H_in[3668])^(data_in[85]&H_in[3669])^(data_in[86]&H_in[3670])^(data_in[87]&H_in[3671])^(data_in[88]&H_in[3672])^(data_in[89]&H_in[3673])^(data_in[90]&H_in[3674])^(data_in[91]&H_in[3675])^(data_in[92]&H_in[3676])^(data_in[93]&H_in[3677])^(data_in[94]&H_in[3678])^(data_in[95]&H_in[3679])^(data_in[96]&H_in[3680])^(data_in[97]&H_in[3681])^(data_in[98]&H_in[3682])^(data_in[99]&H_in[3683])^(data_in[100]&H_in[3684])^(data_in[101]&H_in[3685])^(data_in[102]&H_in[3686])^(data_in[103]&H_in[3687])^(data_in[104]&H_in[3688])^(data_in[105]&H_in[3689])^(data_in[106]&H_in[3690])^(data_in[107]&H_in[3691])^(data_in[108]&H_in[3692])^(data_in[109]&H_in[3693])^(data_in[110]&H_in[3694])^(data_in[111]&H_in[3695])^(data_in[112]&H_in[3696])^(data_in[113]&H_in[3697])^(data_in[114]&H_in[3698])^(data_in[115]&H_in[3699])^(data_in[116]&H_in[3700])^(data_in[117]&H_in[3701])^(data_in[118]&H_in[3702])^(data_in[119]&H_in[3703])^(data_in[120]&H_in[3704])^(data_in[121]&H_in[3705])^(data_in[122]&H_in[3706])^(data_in[123]&H_in[3707])^(data_in[124]&H_in[3708])^(data_in[125]&H_in[3709])^(data_in[126]&H_in[3710])^(data_in[127]&H_in[3711])^(data_in[128]&H_in[3712])^(data_in[129]&H_in[3713])^(data_in[130]&H_in[3714])^(data_in[131]&H_in[3715])^(data_in[132]&H_in[3716])^(data_in[133]&H_in[3717])^(data_in[134]&H_in[3718])^(data_in[135]&H_in[3719])^(data_in[136]&H_in[3720])^(data_in[137]&H_in[3721])^(data_in[138]&H_in[3722])^(data_in[139]&H_in[3723])^(data_in[140]&H_in[3724])^(data_in[141]&H_in[3725])^(data_in[142]&H_in[3726])^(data_in[143]&H_in[3727])^(data_in[144]&H_in[3728])^(data_in[145]&H_in[3729])^(data_in[146]&H_in[3730])^(data_in[147]&H_in[3731])^(data_in[148]&H_in[3732])^(data_in[149]&H_in[3733])^(data_in[150]&H_in[3734])^(data_in[151]&H_in[3735])^(data_in[152]&H_in[3736])^(data_in[153]&H_in[3737])^(data_in[154]&H_in[3738])^(data_in[155]&H_in[3739])^(data_in[156]&H_in[3740])^(data_in[157]&H_in[3741])^(data_in[158]&H_in[3742])^(data_in[159]&H_in[3743])^(data_in[160]&H_in[3744])^(data_in[161]&H_in[3745])^(data_in[162]&H_in[3746])^(data_in[163]&H_in[3747])^(data_in[164]&H_in[3748])^(data_in[165]&H_in[3749])^(data_in[166]&H_in[3750])^(data_in[167]&H_in[3751])^(data_in[168]&H_in[3752])^(data_in[169]&H_in[3753])^(data_in[170]&H_in[3754])^(data_in[171]&H_in[3755])^(data_in[172]&H_in[3756])^(data_in[173]&H_in[3757])^(data_in[174]&H_in[3758])^(data_in[175]&H_in[3759])^(data_in[176]&H_in[3760])^(data_in[177]&H_in[3761])^(data_in[178]&H_in[3762])^(data_in[179]&H_in[3763])^(data_in[180]&H_in[3764])^(data_in[181]&H_in[3765])^(data_in[182]&H_in[3766])^(data_in[183]&H_in[3767])^(data_in[184]&H_in[3768])^(data_in[185]&H_in[3769])^(data_in[186]&H_in[3770])^(data_in[187]&H_in[3771])^(data_in[188]&H_in[3772])^(data_in[189]&H_in[3773])^(data_in[190]&H_in[3774])^(data_in[191]&H_in[3775])^(data_in[192]&H_in[3776])^(data_in[193]&H_in[3777])^(data_in[194]&H_in[3778])^(data_in[195]&H_in[3779])^(data_in[196]&H_in[3780])^(data_in[197]&H_in[3781])^(data_in[198]&H_in[3782])^(data_in[199]&H_in[3783])^(data_in[200]&H_in[3784])^(data_in[201]&H_in[3785])^(data_in[202]&H_in[3786])^(data_in[203]&H_in[3787])^(data_in[204]&H_in[3788])^(data_in[205]&H_in[3789])^(data_in[206]&H_in[3790])^(data_in[207]&H_in[3791])^(data_in[208]&H_in[3792])^(data_in[209]&H_in[3793])^(data_in[210]&H_in[3794])^(data_in[211]&H_in[3795])^(data_in[212]&H_in[3796])^(data_in[213]&H_in[3797])^(data_in[214]&H_in[3798])^(data_in[215]&H_in[3799])^(data_in[216]&H_in[3800])^(data_in[217]&H_in[3801])^(data_in[218]&H_in[3802])^(data_in[219]&H_in[3803])^(data_in[220]&H_in[3804])^(data_in[221]&H_in[3805])^(data_in[222]&H_in[3806])^(data_in[223]&H_in[3807])^(data_in[224]&H_in[3808])^(data_in[225]&H_in[3809])^(data_in[226]&H_in[3810])^(data_in[227]&H_in[3811])^(data_in[228]&H_in[3812])^(data_in[229]&H_in[3813])^(data_in[230]&H_in[3814])^(data_in[231]&H_in[3815])^(data_in[232]&H_in[3816])^(data_in[233]&H_in[3817])^(data_in[234]&H_in[3818])^(data_in[235]&H_in[3819])^(data_in[236]&H_in[3820])^(data_in[237]&H_in[3821])^(data_in[238]&H_in[3822])^(data_in[239]&H_in[3823])^(data_in[240]&H_in[3824])^(data_in[241]&H_in[3825])^(data_in[242]&H_in[3826])^(data_in[243]&H_in[3827])^(data_in[244]&H_in[3828])^(data_in[245]&H_in[3829])^(data_in[246]&H_in[3830])^(data_in[247]&H_in[3831])^(data_in[248]&H_in[3832])^(data_in[249]&H_in[3833])^(data_in[250]&H_in[3834])^(data_in[251]&H_in[3835])^(data_in[252]&H_in[3836])^(data_in[253]&H_in[3837])^(data_in[254]&H_in[3838])^(data_in[255]&H_in[3839]);
         data_out[15]<=(data_in[0]&H_in[3840])^(data_in[1]&H_in[3841])^(data_in[2]&H_in[3842])^(data_in[3]&H_in[3843])^(data_in[4]&H_in[3844])^(data_in[5]&H_in[3845])^(data_in[6]&H_in[3846])^(data_in[7]&H_in[3847])^(data_in[8]&H_in[3848])^(data_in[9]&H_in[3849])^(data_in[10]&H_in[3850])^(data_in[11]&H_in[3851])^(data_in[12]&H_in[3852])^(data_in[13]&H_in[3853])^(data_in[14]&H_in[3854])^(data_in[15]&H_in[3855])^(data_in[16]&H_in[3856])^(data_in[17]&H_in[3857])^(data_in[18]&H_in[3858])^(data_in[19]&H_in[3859])^(data_in[20]&H_in[3860])^(data_in[21]&H_in[3861])^(data_in[22]&H_in[3862])^(data_in[23]&H_in[3863])^(data_in[24]&H_in[3864])^(data_in[25]&H_in[3865])^(data_in[26]&H_in[3866])^(data_in[27]&H_in[3867])^(data_in[28]&H_in[3868])^(data_in[29]&H_in[3869])^(data_in[30]&H_in[3870])^(data_in[31]&H_in[3871])^(data_in[32]&H_in[3872])^(data_in[33]&H_in[3873])^(data_in[34]&H_in[3874])^(data_in[35]&H_in[3875])^(data_in[36]&H_in[3876])^(data_in[37]&H_in[3877])^(data_in[38]&H_in[3878])^(data_in[39]&H_in[3879])^(data_in[40]&H_in[3880])^(data_in[41]&H_in[3881])^(data_in[42]&H_in[3882])^(data_in[43]&H_in[3883])^(data_in[44]&H_in[3884])^(data_in[45]&H_in[3885])^(data_in[46]&H_in[3886])^(data_in[47]&H_in[3887])^(data_in[48]&H_in[3888])^(data_in[49]&H_in[3889])^(data_in[50]&H_in[3890])^(data_in[51]&H_in[3891])^(data_in[52]&H_in[3892])^(data_in[53]&H_in[3893])^(data_in[54]&H_in[3894])^(data_in[55]&H_in[3895])^(data_in[56]&H_in[3896])^(data_in[57]&H_in[3897])^(data_in[58]&H_in[3898])^(data_in[59]&H_in[3899])^(data_in[60]&H_in[3900])^(data_in[61]&H_in[3901])^(data_in[62]&H_in[3902])^(data_in[63]&H_in[3903])^(data_in[64]&H_in[3904])^(data_in[65]&H_in[3905])^(data_in[66]&H_in[3906])^(data_in[67]&H_in[3907])^(data_in[68]&H_in[3908])^(data_in[69]&H_in[3909])^(data_in[70]&H_in[3910])^(data_in[71]&H_in[3911])^(data_in[72]&H_in[3912])^(data_in[73]&H_in[3913])^(data_in[74]&H_in[3914])^(data_in[75]&H_in[3915])^(data_in[76]&H_in[3916])^(data_in[77]&H_in[3917])^(data_in[78]&H_in[3918])^(data_in[79]&H_in[3919])^(data_in[80]&H_in[3920])^(data_in[81]&H_in[3921])^(data_in[82]&H_in[3922])^(data_in[83]&H_in[3923])^(data_in[84]&H_in[3924])^(data_in[85]&H_in[3925])^(data_in[86]&H_in[3926])^(data_in[87]&H_in[3927])^(data_in[88]&H_in[3928])^(data_in[89]&H_in[3929])^(data_in[90]&H_in[3930])^(data_in[91]&H_in[3931])^(data_in[92]&H_in[3932])^(data_in[93]&H_in[3933])^(data_in[94]&H_in[3934])^(data_in[95]&H_in[3935])^(data_in[96]&H_in[3936])^(data_in[97]&H_in[3937])^(data_in[98]&H_in[3938])^(data_in[99]&H_in[3939])^(data_in[100]&H_in[3940])^(data_in[101]&H_in[3941])^(data_in[102]&H_in[3942])^(data_in[103]&H_in[3943])^(data_in[104]&H_in[3944])^(data_in[105]&H_in[3945])^(data_in[106]&H_in[3946])^(data_in[107]&H_in[3947])^(data_in[108]&H_in[3948])^(data_in[109]&H_in[3949])^(data_in[110]&H_in[3950])^(data_in[111]&H_in[3951])^(data_in[112]&H_in[3952])^(data_in[113]&H_in[3953])^(data_in[114]&H_in[3954])^(data_in[115]&H_in[3955])^(data_in[116]&H_in[3956])^(data_in[117]&H_in[3957])^(data_in[118]&H_in[3958])^(data_in[119]&H_in[3959])^(data_in[120]&H_in[3960])^(data_in[121]&H_in[3961])^(data_in[122]&H_in[3962])^(data_in[123]&H_in[3963])^(data_in[124]&H_in[3964])^(data_in[125]&H_in[3965])^(data_in[126]&H_in[3966])^(data_in[127]&H_in[3967])^(data_in[128]&H_in[3968])^(data_in[129]&H_in[3969])^(data_in[130]&H_in[3970])^(data_in[131]&H_in[3971])^(data_in[132]&H_in[3972])^(data_in[133]&H_in[3973])^(data_in[134]&H_in[3974])^(data_in[135]&H_in[3975])^(data_in[136]&H_in[3976])^(data_in[137]&H_in[3977])^(data_in[138]&H_in[3978])^(data_in[139]&H_in[3979])^(data_in[140]&H_in[3980])^(data_in[141]&H_in[3981])^(data_in[142]&H_in[3982])^(data_in[143]&H_in[3983])^(data_in[144]&H_in[3984])^(data_in[145]&H_in[3985])^(data_in[146]&H_in[3986])^(data_in[147]&H_in[3987])^(data_in[148]&H_in[3988])^(data_in[149]&H_in[3989])^(data_in[150]&H_in[3990])^(data_in[151]&H_in[3991])^(data_in[152]&H_in[3992])^(data_in[153]&H_in[3993])^(data_in[154]&H_in[3994])^(data_in[155]&H_in[3995])^(data_in[156]&H_in[3996])^(data_in[157]&H_in[3997])^(data_in[158]&H_in[3998])^(data_in[159]&H_in[3999])^(data_in[160]&H_in[4000])^(data_in[161]&H_in[4001])^(data_in[162]&H_in[4002])^(data_in[163]&H_in[4003])^(data_in[164]&H_in[4004])^(data_in[165]&H_in[4005])^(data_in[166]&H_in[4006])^(data_in[167]&H_in[4007])^(data_in[168]&H_in[4008])^(data_in[169]&H_in[4009])^(data_in[170]&H_in[4010])^(data_in[171]&H_in[4011])^(data_in[172]&H_in[4012])^(data_in[173]&H_in[4013])^(data_in[174]&H_in[4014])^(data_in[175]&H_in[4015])^(data_in[176]&H_in[4016])^(data_in[177]&H_in[4017])^(data_in[178]&H_in[4018])^(data_in[179]&H_in[4019])^(data_in[180]&H_in[4020])^(data_in[181]&H_in[4021])^(data_in[182]&H_in[4022])^(data_in[183]&H_in[4023])^(data_in[184]&H_in[4024])^(data_in[185]&H_in[4025])^(data_in[186]&H_in[4026])^(data_in[187]&H_in[4027])^(data_in[188]&H_in[4028])^(data_in[189]&H_in[4029])^(data_in[190]&H_in[4030])^(data_in[191]&H_in[4031])^(data_in[192]&H_in[4032])^(data_in[193]&H_in[4033])^(data_in[194]&H_in[4034])^(data_in[195]&H_in[4035])^(data_in[196]&H_in[4036])^(data_in[197]&H_in[4037])^(data_in[198]&H_in[4038])^(data_in[199]&H_in[4039])^(data_in[200]&H_in[4040])^(data_in[201]&H_in[4041])^(data_in[202]&H_in[4042])^(data_in[203]&H_in[4043])^(data_in[204]&H_in[4044])^(data_in[205]&H_in[4045])^(data_in[206]&H_in[4046])^(data_in[207]&H_in[4047])^(data_in[208]&H_in[4048])^(data_in[209]&H_in[4049])^(data_in[210]&H_in[4050])^(data_in[211]&H_in[4051])^(data_in[212]&H_in[4052])^(data_in[213]&H_in[4053])^(data_in[214]&H_in[4054])^(data_in[215]&H_in[4055])^(data_in[216]&H_in[4056])^(data_in[217]&H_in[4057])^(data_in[218]&H_in[4058])^(data_in[219]&H_in[4059])^(data_in[220]&H_in[4060])^(data_in[221]&H_in[4061])^(data_in[222]&H_in[4062])^(data_in[223]&H_in[4063])^(data_in[224]&H_in[4064])^(data_in[225]&H_in[4065])^(data_in[226]&H_in[4066])^(data_in[227]&H_in[4067])^(data_in[228]&H_in[4068])^(data_in[229]&H_in[4069])^(data_in[230]&H_in[4070])^(data_in[231]&H_in[4071])^(data_in[232]&H_in[4072])^(data_in[233]&H_in[4073])^(data_in[234]&H_in[4074])^(data_in[235]&H_in[4075])^(data_in[236]&H_in[4076])^(data_in[237]&H_in[4077])^(data_in[238]&H_in[4078])^(data_in[239]&H_in[4079])^(data_in[240]&H_in[4080])^(data_in[241]&H_in[4081])^(data_in[242]&H_in[4082])^(data_in[243]&H_in[4083])^(data_in[244]&H_in[4084])^(data_in[245]&H_in[4085])^(data_in[246]&H_in[4086])^(data_in[247]&H_in[4087])^(data_in[248]&H_in[4088])^(data_in[249]&H_in[4089])^(data_in[250]&H_in[4090])^(data_in[251]&H_in[4091])^(data_in[252]&H_in[4092])^(data_in[253]&H_in[4093])^(data_in[254]&H_in[4094])^(data_in[255]&H_in[4095]);
          
         end
         else if(r_en==0&&cnt==1)begin
         data_out[0]<=data_out[0]^(data_in[0]&H_in[0])^(data_in[1]&H_in[1])^(data_in[2]&H_in[2])^(data_in[3]&H_in[3])^(data_in[4]&H_in[4])^(data_in[5]&H_in[5])^(data_in[6]&H_in[6])^(data_in[7]&H_in[7])^(data_in[8]&H_in[8])^(data_in[9]&H_in[9])^(data_in[10]&H_in[10])^(data_in[11]&H_in[11])^(data_in[12]&H_in[12])^(data_in[13]&H_in[13])^(data_in[14]&H_in[14])^(data_in[15]&H_in[15])^(data_in[16]&H_in[16])^(data_in[17]&H_in[17])^(data_in[18]&H_in[18])^(data_in[19]&H_in[19])^(data_in[20]&H_in[20])^(data_in[21]&H_in[21])^(data_in[22]&H_in[22])^(data_in[23]&H_in[23])^(data_in[24]&H_in[24])^(data_in[25]&H_in[25])^(data_in[26]&H_in[26])^(data_in[27]&H_in[27])^(data_in[28]&H_in[28])^(data_in[29]&H_in[29])^(data_in[30]&H_in[30])^(data_in[31]&H_in[31])^(data_in[32]&H_in[32])^(data_in[33]&H_in[33])^(data_in[34]&H_in[34])^(data_in[35]&H_in[35])^(data_in[36]&H_in[36])^(data_in[37]&H_in[37])^(data_in[38]&H_in[38])^(data_in[39]&H_in[39])^(data_in[40]&H_in[40])^(data_in[41]&H_in[41])^(data_in[42]&H_in[42])^(data_in[43]&H_in[43])^(data_in[44]&H_in[44])^(data_in[45]&H_in[45])^(data_in[46]&H_in[46])^(data_in[47]&H_in[47])^(data_in[48]&H_in[48])^(data_in[49]&H_in[49])^(data_in[50]&H_in[50])^(data_in[51]&H_in[51])^(data_in[52]&H_in[52])^(data_in[53]&H_in[53])^(data_in[54]&H_in[54])^(data_in[55]&H_in[55])^(data_in[56]&H_in[56])^(data_in[57]&H_in[57])^(data_in[58]&H_in[58])^(data_in[59]&H_in[59])^(data_in[60]&H_in[60])^(data_in[61]&H_in[61])^(data_in[62]&H_in[62])^(data_in[63]&H_in[63])^(data_in[64]&H_in[64])^(data_in[65]&H_in[65])^(data_in[66]&H_in[66])^(data_in[67]&H_in[67])^(data_in[68]&H_in[68])^(data_in[69]&H_in[69])^(data_in[70]&H_in[70])^(data_in[71]&H_in[71])^(data_in[72]&H_in[72])^(data_in[73]&H_in[73])^(data_in[74]&H_in[74])^(data_in[75]&H_in[75])^(data_in[76]&H_in[76])^(data_in[77]&H_in[77])^(data_in[78]&H_in[78])^(data_in[79]&H_in[79])^(data_in[80]&H_in[80])^(data_in[81]&H_in[81])^(data_in[82]&H_in[82])^(data_in[83]&H_in[83])^(data_in[84]&H_in[84])^(data_in[85]&H_in[85])^(data_in[86]&H_in[86])^(data_in[87]&H_in[87])^(data_in[88]&H_in[88])^(data_in[89]&H_in[89])^(data_in[90]&H_in[90])^(data_in[91]&H_in[91])^(data_in[92]&H_in[92])^(data_in[93]&H_in[93])^(data_in[94]&H_in[94])^(data_in[95]&H_in[95])^(data_in[96]&H_in[96])^(data_in[97]&H_in[97])^(data_in[98]&H_in[98])^(data_in[99]&H_in[99])^(data_in[100]&H_in[100])^(data_in[101]&H_in[101])^(data_in[102]&H_in[102])^(data_in[103]&H_in[103])^(data_in[104]&H_in[104])^(data_in[105]&H_in[105])^(data_in[106]&H_in[106])^(data_in[107]&H_in[107])^(data_in[108]&H_in[108])^(data_in[109]&H_in[109])^(data_in[110]&H_in[110])^(data_in[111]&H_in[111])^(data_in[112]&H_in[112])^(data_in[113]&H_in[113])^(data_in[114]&H_in[114])^(data_in[115]&H_in[115])^(data_in[116]&H_in[116])^(data_in[117]&H_in[117])^(data_in[118]&H_in[118])^(data_in[119]&H_in[119])^(data_in[120]&H_in[120])^(data_in[121]&H_in[121])^(data_in[122]&H_in[122])^(data_in[123]&H_in[123])^(data_in[124]&H_in[124])^(data_in[125]&H_in[125])^(data_in[126]&H_in[126])^(data_in[127]&H_in[127])^(data_in[128]&H_in[128])^(data_in[129]&H_in[129])^(data_in[130]&H_in[130])^(data_in[131]&H_in[131])^(data_in[132]&H_in[132])^(data_in[133]&H_in[133])^(data_in[134]&H_in[134])^(data_in[135]&H_in[135])^(data_in[136]&H_in[136])^(data_in[137]&H_in[137])^(data_in[138]&H_in[138])^(data_in[139]&H_in[139])^(data_in[140]&H_in[140])^(data_in[141]&H_in[141])^(data_in[142]&H_in[142])^(data_in[143]&H_in[143])^(data_in[144]&H_in[144])^(data_in[145]&H_in[145])^(data_in[146]&H_in[146])^(data_in[147]&H_in[147])^(data_in[148]&H_in[148])^(data_in[149]&H_in[149])^(data_in[150]&H_in[150])^(data_in[151]&H_in[151])^(data_in[152]&H_in[152])^(data_in[153]&H_in[153])^(data_in[154]&H_in[154])^(data_in[155]&H_in[155])^(data_in[156]&H_in[156])^(data_in[157]&H_in[157])^(data_in[158]&H_in[158])^(data_in[159]&H_in[159])^(data_in[160]&H_in[160])^(data_in[161]&H_in[161])^(data_in[162]&H_in[162])^(data_in[163]&H_in[163])^(data_in[164]&H_in[164])^(data_in[165]&H_in[165])^(data_in[166]&H_in[166])^(data_in[167]&H_in[167])^(data_in[168]&H_in[168])^(data_in[169]&H_in[169])^(data_in[170]&H_in[170])^(data_in[171]&H_in[171])^(data_in[172]&H_in[172])^(data_in[173]&H_in[173])^(data_in[174]&H_in[174])^(data_in[175]&H_in[175])^(data_in[176]&H_in[176])^(data_in[177]&H_in[177])^(data_in[178]&H_in[178])^(data_in[179]&H_in[179])^(data_in[180]&H_in[180])^(data_in[181]&H_in[181])^(data_in[182]&H_in[182])^(data_in[183]&H_in[183])^(data_in[184]&H_in[184])^(data_in[185]&H_in[185])^(data_in[186]&H_in[186])^(data_in[187]&H_in[187])^(data_in[188]&H_in[188])^(data_in[189]&H_in[189])^(data_in[190]&H_in[190])^(data_in[191]&H_in[191])^(data_in[192]&H_in[192])^(data_in[193]&H_in[193])^(data_in[194]&H_in[194])^(data_in[195]&H_in[195])^(data_in[196]&H_in[196])^(data_in[197]&H_in[197])^(data_in[198]&H_in[198])^(data_in[199]&H_in[199])^(data_in[200]&H_in[200])^(data_in[201]&H_in[201])^(data_in[202]&H_in[202])^(data_in[203]&H_in[203])^(data_in[204]&H_in[204])^(data_in[205]&H_in[205])^(data_in[206]&H_in[206])^(data_in[207]&H_in[207])^(data_in[208]&H_in[208])^(data_in[209]&H_in[209])^(data_in[210]&H_in[210])^(data_in[211]&H_in[211])^(data_in[212]&H_in[212])^(data_in[213]&H_in[213])^(data_in[214]&H_in[214])^(data_in[215]&H_in[215])^(data_in[216]&H_in[216])^(data_in[217]&H_in[217])^(data_in[218]&H_in[218])^(data_in[219]&H_in[219])^(data_in[220]&H_in[220])^(data_in[221]&H_in[221])^(data_in[222]&H_in[222])^(data_in[223]&H_in[223])^(data_in[224]&H_in[224])^(data_in[225]&H_in[225])^(data_in[226]&H_in[226])^(data_in[227]&H_in[227])^(data_in[228]&H_in[228])^(data_in[229]&H_in[229])^(data_in[230]&H_in[230])^(data_in[231]&H_in[231])^(data_in[232]&H_in[232])^(data_in[233]&H_in[233])^(data_in[234]&H_in[234])^(data_in[235]&H_in[235])^(data_in[236]&H_in[236])^(data_in[237]&H_in[237])^(data_in[238]&H_in[238])^(data_in[239]&H_in[239])^(data_in[240]&H_in[240])^(data_in[241]&H_in[241])^(data_in[242]&H_in[242])^(data_in[243]&H_in[243])^(data_in[244]&H_in[244])^(data_in[245]&H_in[245])^(data_in[246]&H_in[246])^(data_in[247]&H_in[247])^(data_in[248]&H_in[248])^(data_in[249]&H_in[249])^(data_in[250]&H_in[250])^(data_in[251]&H_in[251])^(data_in[252]&H_in[252])^(data_in[253]&H_in[253])^(data_in[254]&H_in[254])^(data_in[255]&H_in[255]);
         data_out[1]<=data_out[1]^(data_in[0]&H_in[256])^(data_in[1]&H_in[257])^(data_in[2]&H_in[258])^(data_in[3]&H_in[259])^(data_in[4]&H_in[260])^(data_in[5]&H_in[261])^(data_in[6]&H_in[262])^(data_in[7]&H_in[263])^(data_in[8]&H_in[264])^(data_in[9]&H_in[265])^(data_in[10]&H_in[266])^(data_in[11]&H_in[267])^(data_in[12]&H_in[268])^(data_in[13]&H_in[269])^(data_in[14]&H_in[270])^(data_in[15]&H_in[271])^(data_in[16]&H_in[272])^(data_in[17]&H_in[273])^(data_in[18]&H_in[274])^(data_in[19]&H_in[275])^(data_in[20]&H_in[276])^(data_in[21]&H_in[277])^(data_in[22]&H_in[278])^(data_in[23]&H_in[279])^(data_in[24]&H_in[280])^(data_in[25]&H_in[281])^(data_in[26]&H_in[282])^(data_in[27]&H_in[283])^(data_in[28]&H_in[284])^(data_in[29]&H_in[285])^(data_in[30]&H_in[286])^(data_in[31]&H_in[287])^(data_in[32]&H_in[288])^(data_in[33]&H_in[289])^(data_in[34]&H_in[290])^(data_in[35]&H_in[291])^(data_in[36]&H_in[292])^(data_in[37]&H_in[293])^(data_in[38]&H_in[294])^(data_in[39]&H_in[295])^(data_in[40]&H_in[296])^(data_in[41]&H_in[297])^(data_in[42]&H_in[298])^(data_in[43]&H_in[299])^(data_in[44]&H_in[300])^(data_in[45]&H_in[301])^(data_in[46]&H_in[302])^(data_in[47]&H_in[303])^(data_in[48]&H_in[304])^(data_in[49]&H_in[305])^(data_in[50]&H_in[306])^(data_in[51]&H_in[307])^(data_in[52]&H_in[308])^(data_in[53]&H_in[309])^(data_in[54]&H_in[310])^(data_in[55]&H_in[311])^(data_in[56]&H_in[312])^(data_in[57]&H_in[313])^(data_in[58]&H_in[314])^(data_in[59]&H_in[315])^(data_in[60]&H_in[316])^(data_in[61]&H_in[317])^(data_in[62]&H_in[318])^(data_in[63]&H_in[319])^(data_in[64]&H_in[320])^(data_in[65]&H_in[321])^(data_in[66]&H_in[322])^(data_in[67]&H_in[323])^(data_in[68]&H_in[324])^(data_in[69]&H_in[325])^(data_in[70]&H_in[326])^(data_in[71]&H_in[327])^(data_in[72]&H_in[328])^(data_in[73]&H_in[329])^(data_in[74]&H_in[330])^(data_in[75]&H_in[331])^(data_in[76]&H_in[332])^(data_in[77]&H_in[333])^(data_in[78]&H_in[334])^(data_in[79]&H_in[335])^(data_in[80]&H_in[336])^(data_in[81]&H_in[337])^(data_in[82]&H_in[338])^(data_in[83]&H_in[339])^(data_in[84]&H_in[340])^(data_in[85]&H_in[341])^(data_in[86]&H_in[342])^(data_in[87]&H_in[343])^(data_in[88]&H_in[344])^(data_in[89]&H_in[345])^(data_in[90]&H_in[346])^(data_in[91]&H_in[347])^(data_in[92]&H_in[348])^(data_in[93]&H_in[349])^(data_in[94]&H_in[350])^(data_in[95]&H_in[351])^(data_in[96]&H_in[352])^(data_in[97]&H_in[353])^(data_in[98]&H_in[354])^(data_in[99]&H_in[355])^(data_in[100]&H_in[356])^(data_in[101]&H_in[357])^(data_in[102]&H_in[358])^(data_in[103]&H_in[359])^(data_in[104]&H_in[360])^(data_in[105]&H_in[361])^(data_in[106]&H_in[362])^(data_in[107]&H_in[363])^(data_in[108]&H_in[364])^(data_in[109]&H_in[365])^(data_in[110]&H_in[366])^(data_in[111]&H_in[367])^(data_in[112]&H_in[368])^(data_in[113]&H_in[369])^(data_in[114]&H_in[370])^(data_in[115]&H_in[371])^(data_in[116]&H_in[372])^(data_in[117]&H_in[373])^(data_in[118]&H_in[374])^(data_in[119]&H_in[375])^(data_in[120]&H_in[376])^(data_in[121]&H_in[377])^(data_in[122]&H_in[378])^(data_in[123]&H_in[379])^(data_in[124]&H_in[380])^(data_in[125]&H_in[381])^(data_in[126]&H_in[382])^(data_in[127]&H_in[383])^(data_in[128]&H_in[384])^(data_in[129]&H_in[385])^(data_in[130]&H_in[386])^(data_in[131]&H_in[387])^(data_in[132]&H_in[388])^(data_in[133]&H_in[389])^(data_in[134]&H_in[390])^(data_in[135]&H_in[391])^(data_in[136]&H_in[392])^(data_in[137]&H_in[393])^(data_in[138]&H_in[394])^(data_in[139]&H_in[395])^(data_in[140]&H_in[396])^(data_in[141]&H_in[397])^(data_in[142]&H_in[398])^(data_in[143]&H_in[399])^(data_in[144]&H_in[400])^(data_in[145]&H_in[401])^(data_in[146]&H_in[402])^(data_in[147]&H_in[403])^(data_in[148]&H_in[404])^(data_in[149]&H_in[405])^(data_in[150]&H_in[406])^(data_in[151]&H_in[407])^(data_in[152]&H_in[408])^(data_in[153]&H_in[409])^(data_in[154]&H_in[410])^(data_in[155]&H_in[411])^(data_in[156]&H_in[412])^(data_in[157]&H_in[413])^(data_in[158]&H_in[414])^(data_in[159]&H_in[415])^(data_in[160]&H_in[416])^(data_in[161]&H_in[417])^(data_in[162]&H_in[418])^(data_in[163]&H_in[419])^(data_in[164]&H_in[420])^(data_in[165]&H_in[421])^(data_in[166]&H_in[422])^(data_in[167]&H_in[423])^(data_in[168]&H_in[424])^(data_in[169]&H_in[425])^(data_in[170]&H_in[426])^(data_in[171]&H_in[427])^(data_in[172]&H_in[428])^(data_in[173]&H_in[429])^(data_in[174]&H_in[430])^(data_in[175]&H_in[431])^(data_in[176]&H_in[432])^(data_in[177]&H_in[433])^(data_in[178]&H_in[434])^(data_in[179]&H_in[435])^(data_in[180]&H_in[436])^(data_in[181]&H_in[437])^(data_in[182]&H_in[438])^(data_in[183]&H_in[439])^(data_in[184]&H_in[440])^(data_in[185]&H_in[441])^(data_in[186]&H_in[442])^(data_in[187]&H_in[443])^(data_in[188]&H_in[444])^(data_in[189]&H_in[445])^(data_in[190]&H_in[446])^(data_in[191]&H_in[447])^(data_in[192]&H_in[448])^(data_in[193]&H_in[449])^(data_in[194]&H_in[450])^(data_in[195]&H_in[451])^(data_in[196]&H_in[452])^(data_in[197]&H_in[453])^(data_in[198]&H_in[454])^(data_in[199]&H_in[455])^(data_in[200]&H_in[456])^(data_in[201]&H_in[457])^(data_in[202]&H_in[458])^(data_in[203]&H_in[459])^(data_in[204]&H_in[460])^(data_in[205]&H_in[461])^(data_in[206]&H_in[462])^(data_in[207]&H_in[463])^(data_in[208]&H_in[464])^(data_in[209]&H_in[465])^(data_in[210]&H_in[466])^(data_in[211]&H_in[467])^(data_in[212]&H_in[468])^(data_in[213]&H_in[469])^(data_in[214]&H_in[470])^(data_in[215]&H_in[471])^(data_in[216]&H_in[472])^(data_in[217]&H_in[473])^(data_in[218]&H_in[474])^(data_in[219]&H_in[475])^(data_in[220]&H_in[476])^(data_in[221]&H_in[477])^(data_in[222]&H_in[478])^(data_in[223]&H_in[479])^(data_in[224]&H_in[480])^(data_in[225]&H_in[481])^(data_in[226]&H_in[482])^(data_in[227]&H_in[483])^(data_in[228]&H_in[484])^(data_in[229]&H_in[485])^(data_in[230]&H_in[486])^(data_in[231]&H_in[487])^(data_in[232]&H_in[488])^(data_in[233]&H_in[489])^(data_in[234]&H_in[490])^(data_in[235]&H_in[491])^(data_in[236]&H_in[492])^(data_in[237]&H_in[493])^(data_in[238]&H_in[494])^(data_in[239]&H_in[495])^(data_in[240]&H_in[496])^(data_in[241]&H_in[497])^(data_in[242]&H_in[498])^(data_in[243]&H_in[499])^(data_in[244]&H_in[500])^(data_in[245]&H_in[501])^(data_in[246]&H_in[502])^(data_in[247]&H_in[503])^(data_in[248]&H_in[504])^(data_in[249]&H_in[505])^(data_in[250]&H_in[506])^(data_in[251]&H_in[507])^(data_in[252]&H_in[508])^(data_in[253]&H_in[509])^(data_in[254]&H_in[510])^(data_in[255]&H_in[511]);
         data_out[2]<=data_out[2]^(data_in[0]&H_in[512])^(data_in[1]&H_in[513])^(data_in[2]&H_in[514])^(data_in[3]&H_in[515])^(data_in[4]&H_in[516])^(data_in[5]&H_in[517])^(data_in[6]&H_in[518])^(data_in[7]&H_in[519])^(data_in[8]&H_in[520])^(data_in[9]&H_in[521])^(data_in[10]&H_in[522])^(data_in[11]&H_in[523])^(data_in[12]&H_in[524])^(data_in[13]&H_in[525])^(data_in[14]&H_in[526])^(data_in[15]&H_in[527])^(data_in[16]&H_in[528])^(data_in[17]&H_in[529])^(data_in[18]&H_in[530])^(data_in[19]&H_in[531])^(data_in[20]&H_in[532])^(data_in[21]&H_in[533])^(data_in[22]&H_in[534])^(data_in[23]&H_in[535])^(data_in[24]&H_in[536])^(data_in[25]&H_in[537])^(data_in[26]&H_in[538])^(data_in[27]&H_in[539])^(data_in[28]&H_in[540])^(data_in[29]&H_in[541])^(data_in[30]&H_in[542])^(data_in[31]&H_in[543])^(data_in[32]&H_in[544])^(data_in[33]&H_in[545])^(data_in[34]&H_in[546])^(data_in[35]&H_in[547])^(data_in[36]&H_in[548])^(data_in[37]&H_in[549])^(data_in[38]&H_in[550])^(data_in[39]&H_in[551])^(data_in[40]&H_in[552])^(data_in[41]&H_in[553])^(data_in[42]&H_in[554])^(data_in[43]&H_in[555])^(data_in[44]&H_in[556])^(data_in[45]&H_in[557])^(data_in[46]&H_in[558])^(data_in[47]&H_in[559])^(data_in[48]&H_in[560])^(data_in[49]&H_in[561])^(data_in[50]&H_in[562])^(data_in[51]&H_in[563])^(data_in[52]&H_in[564])^(data_in[53]&H_in[565])^(data_in[54]&H_in[566])^(data_in[55]&H_in[567])^(data_in[56]&H_in[568])^(data_in[57]&H_in[569])^(data_in[58]&H_in[570])^(data_in[59]&H_in[571])^(data_in[60]&H_in[572])^(data_in[61]&H_in[573])^(data_in[62]&H_in[574])^(data_in[63]&H_in[575])^(data_in[64]&H_in[576])^(data_in[65]&H_in[577])^(data_in[66]&H_in[578])^(data_in[67]&H_in[579])^(data_in[68]&H_in[580])^(data_in[69]&H_in[581])^(data_in[70]&H_in[582])^(data_in[71]&H_in[583])^(data_in[72]&H_in[584])^(data_in[73]&H_in[585])^(data_in[74]&H_in[586])^(data_in[75]&H_in[587])^(data_in[76]&H_in[588])^(data_in[77]&H_in[589])^(data_in[78]&H_in[590])^(data_in[79]&H_in[591])^(data_in[80]&H_in[592])^(data_in[81]&H_in[593])^(data_in[82]&H_in[594])^(data_in[83]&H_in[595])^(data_in[84]&H_in[596])^(data_in[85]&H_in[597])^(data_in[86]&H_in[598])^(data_in[87]&H_in[599])^(data_in[88]&H_in[600])^(data_in[89]&H_in[601])^(data_in[90]&H_in[602])^(data_in[91]&H_in[603])^(data_in[92]&H_in[604])^(data_in[93]&H_in[605])^(data_in[94]&H_in[606])^(data_in[95]&H_in[607])^(data_in[96]&H_in[608])^(data_in[97]&H_in[609])^(data_in[98]&H_in[610])^(data_in[99]&H_in[611])^(data_in[100]&H_in[612])^(data_in[101]&H_in[613])^(data_in[102]&H_in[614])^(data_in[103]&H_in[615])^(data_in[104]&H_in[616])^(data_in[105]&H_in[617])^(data_in[106]&H_in[618])^(data_in[107]&H_in[619])^(data_in[108]&H_in[620])^(data_in[109]&H_in[621])^(data_in[110]&H_in[622])^(data_in[111]&H_in[623])^(data_in[112]&H_in[624])^(data_in[113]&H_in[625])^(data_in[114]&H_in[626])^(data_in[115]&H_in[627])^(data_in[116]&H_in[628])^(data_in[117]&H_in[629])^(data_in[118]&H_in[630])^(data_in[119]&H_in[631])^(data_in[120]&H_in[632])^(data_in[121]&H_in[633])^(data_in[122]&H_in[634])^(data_in[123]&H_in[635])^(data_in[124]&H_in[636])^(data_in[125]&H_in[637])^(data_in[126]&H_in[638])^(data_in[127]&H_in[639])^(data_in[128]&H_in[640])^(data_in[129]&H_in[641])^(data_in[130]&H_in[642])^(data_in[131]&H_in[643])^(data_in[132]&H_in[644])^(data_in[133]&H_in[645])^(data_in[134]&H_in[646])^(data_in[135]&H_in[647])^(data_in[136]&H_in[648])^(data_in[137]&H_in[649])^(data_in[138]&H_in[650])^(data_in[139]&H_in[651])^(data_in[140]&H_in[652])^(data_in[141]&H_in[653])^(data_in[142]&H_in[654])^(data_in[143]&H_in[655])^(data_in[144]&H_in[656])^(data_in[145]&H_in[657])^(data_in[146]&H_in[658])^(data_in[147]&H_in[659])^(data_in[148]&H_in[660])^(data_in[149]&H_in[661])^(data_in[150]&H_in[662])^(data_in[151]&H_in[663])^(data_in[152]&H_in[664])^(data_in[153]&H_in[665])^(data_in[154]&H_in[666])^(data_in[155]&H_in[667])^(data_in[156]&H_in[668])^(data_in[157]&H_in[669])^(data_in[158]&H_in[670])^(data_in[159]&H_in[671])^(data_in[160]&H_in[672])^(data_in[161]&H_in[673])^(data_in[162]&H_in[674])^(data_in[163]&H_in[675])^(data_in[164]&H_in[676])^(data_in[165]&H_in[677])^(data_in[166]&H_in[678])^(data_in[167]&H_in[679])^(data_in[168]&H_in[680])^(data_in[169]&H_in[681])^(data_in[170]&H_in[682])^(data_in[171]&H_in[683])^(data_in[172]&H_in[684])^(data_in[173]&H_in[685])^(data_in[174]&H_in[686])^(data_in[175]&H_in[687])^(data_in[176]&H_in[688])^(data_in[177]&H_in[689])^(data_in[178]&H_in[690])^(data_in[179]&H_in[691])^(data_in[180]&H_in[692])^(data_in[181]&H_in[693])^(data_in[182]&H_in[694])^(data_in[183]&H_in[695])^(data_in[184]&H_in[696])^(data_in[185]&H_in[697])^(data_in[186]&H_in[698])^(data_in[187]&H_in[699])^(data_in[188]&H_in[700])^(data_in[189]&H_in[701])^(data_in[190]&H_in[702])^(data_in[191]&H_in[703])^(data_in[192]&H_in[704])^(data_in[193]&H_in[705])^(data_in[194]&H_in[706])^(data_in[195]&H_in[707])^(data_in[196]&H_in[708])^(data_in[197]&H_in[709])^(data_in[198]&H_in[710])^(data_in[199]&H_in[711])^(data_in[200]&H_in[712])^(data_in[201]&H_in[713])^(data_in[202]&H_in[714])^(data_in[203]&H_in[715])^(data_in[204]&H_in[716])^(data_in[205]&H_in[717])^(data_in[206]&H_in[718])^(data_in[207]&H_in[719])^(data_in[208]&H_in[720])^(data_in[209]&H_in[721])^(data_in[210]&H_in[722])^(data_in[211]&H_in[723])^(data_in[212]&H_in[724])^(data_in[213]&H_in[725])^(data_in[214]&H_in[726])^(data_in[215]&H_in[727])^(data_in[216]&H_in[728])^(data_in[217]&H_in[729])^(data_in[218]&H_in[730])^(data_in[219]&H_in[731])^(data_in[220]&H_in[732])^(data_in[221]&H_in[733])^(data_in[222]&H_in[734])^(data_in[223]&H_in[735])^(data_in[224]&H_in[736])^(data_in[225]&H_in[737])^(data_in[226]&H_in[738])^(data_in[227]&H_in[739])^(data_in[228]&H_in[740])^(data_in[229]&H_in[741])^(data_in[230]&H_in[742])^(data_in[231]&H_in[743])^(data_in[232]&H_in[744])^(data_in[233]&H_in[745])^(data_in[234]&H_in[746])^(data_in[235]&H_in[747])^(data_in[236]&H_in[748])^(data_in[237]&H_in[749])^(data_in[238]&H_in[750])^(data_in[239]&H_in[751])^(data_in[240]&H_in[752])^(data_in[241]&H_in[753])^(data_in[242]&H_in[754])^(data_in[243]&H_in[755])^(data_in[244]&H_in[756])^(data_in[245]&H_in[757])^(data_in[246]&H_in[758])^(data_in[247]&H_in[759])^(data_in[248]&H_in[760])^(data_in[249]&H_in[761])^(data_in[250]&H_in[762])^(data_in[251]&H_in[763])^(data_in[252]&H_in[764])^(data_in[253]&H_in[765])^(data_in[254]&H_in[766])^(data_in[255]&H_in[767]);
         data_out[3]<=data_out[3]^(data_in[0]&H_in[768])^(data_in[1]&H_in[769])^(data_in[2]&H_in[770])^(data_in[3]&H_in[771])^(data_in[4]&H_in[772])^(data_in[5]&H_in[773])^(data_in[6]&H_in[774])^(data_in[7]&H_in[775])^(data_in[8]&H_in[776])^(data_in[9]&H_in[777])^(data_in[10]&H_in[778])^(data_in[11]&H_in[779])^(data_in[12]&H_in[780])^(data_in[13]&H_in[781])^(data_in[14]&H_in[782])^(data_in[15]&H_in[783])^(data_in[16]&H_in[784])^(data_in[17]&H_in[785])^(data_in[18]&H_in[786])^(data_in[19]&H_in[787])^(data_in[20]&H_in[788])^(data_in[21]&H_in[789])^(data_in[22]&H_in[790])^(data_in[23]&H_in[791])^(data_in[24]&H_in[792])^(data_in[25]&H_in[793])^(data_in[26]&H_in[794])^(data_in[27]&H_in[795])^(data_in[28]&H_in[796])^(data_in[29]&H_in[797])^(data_in[30]&H_in[798])^(data_in[31]&H_in[799])^(data_in[32]&H_in[800])^(data_in[33]&H_in[801])^(data_in[34]&H_in[802])^(data_in[35]&H_in[803])^(data_in[36]&H_in[804])^(data_in[37]&H_in[805])^(data_in[38]&H_in[806])^(data_in[39]&H_in[807])^(data_in[40]&H_in[808])^(data_in[41]&H_in[809])^(data_in[42]&H_in[810])^(data_in[43]&H_in[811])^(data_in[44]&H_in[812])^(data_in[45]&H_in[813])^(data_in[46]&H_in[814])^(data_in[47]&H_in[815])^(data_in[48]&H_in[816])^(data_in[49]&H_in[817])^(data_in[50]&H_in[818])^(data_in[51]&H_in[819])^(data_in[52]&H_in[820])^(data_in[53]&H_in[821])^(data_in[54]&H_in[822])^(data_in[55]&H_in[823])^(data_in[56]&H_in[824])^(data_in[57]&H_in[825])^(data_in[58]&H_in[826])^(data_in[59]&H_in[827])^(data_in[60]&H_in[828])^(data_in[61]&H_in[829])^(data_in[62]&H_in[830])^(data_in[63]&H_in[831])^(data_in[64]&H_in[832])^(data_in[65]&H_in[833])^(data_in[66]&H_in[834])^(data_in[67]&H_in[835])^(data_in[68]&H_in[836])^(data_in[69]&H_in[837])^(data_in[70]&H_in[838])^(data_in[71]&H_in[839])^(data_in[72]&H_in[840])^(data_in[73]&H_in[841])^(data_in[74]&H_in[842])^(data_in[75]&H_in[843])^(data_in[76]&H_in[844])^(data_in[77]&H_in[845])^(data_in[78]&H_in[846])^(data_in[79]&H_in[847])^(data_in[80]&H_in[848])^(data_in[81]&H_in[849])^(data_in[82]&H_in[850])^(data_in[83]&H_in[851])^(data_in[84]&H_in[852])^(data_in[85]&H_in[853])^(data_in[86]&H_in[854])^(data_in[87]&H_in[855])^(data_in[88]&H_in[856])^(data_in[89]&H_in[857])^(data_in[90]&H_in[858])^(data_in[91]&H_in[859])^(data_in[92]&H_in[860])^(data_in[93]&H_in[861])^(data_in[94]&H_in[862])^(data_in[95]&H_in[863])^(data_in[96]&H_in[864])^(data_in[97]&H_in[865])^(data_in[98]&H_in[866])^(data_in[99]&H_in[867])^(data_in[100]&H_in[868])^(data_in[101]&H_in[869])^(data_in[102]&H_in[870])^(data_in[103]&H_in[871])^(data_in[104]&H_in[872])^(data_in[105]&H_in[873])^(data_in[106]&H_in[874])^(data_in[107]&H_in[875])^(data_in[108]&H_in[876])^(data_in[109]&H_in[877])^(data_in[110]&H_in[878])^(data_in[111]&H_in[879])^(data_in[112]&H_in[880])^(data_in[113]&H_in[881])^(data_in[114]&H_in[882])^(data_in[115]&H_in[883])^(data_in[116]&H_in[884])^(data_in[117]&H_in[885])^(data_in[118]&H_in[886])^(data_in[119]&H_in[887])^(data_in[120]&H_in[888])^(data_in[121]&H_in[889])^(data_in[122]&H_in[890])^(data_in[123]&H_in[891])^(data_in[124]&H_in[892])^(data_in[125]&H_in[893])^(data_in[126]&H_in[894])^(data_in[127]&H_in[895])^(data_in[128]&H_in[896])^(data_in[129]&H_in[897])^(data_in[130]&H_in[898])^(data_in[131]&H_in[899])^(data_in[132]&H_in[900])^(data_in[133]&H_in[901])^(data_in[134]&H_in[902])^(data_in[135]&H_in[903])^(data_in[136]&H_in[904])^(data_in[137]&H_in[905])^(data_in[138]&H_in[906])^(data_in[139]&H_in[907])^(data_in[140]&H_in[908])^(data_in[141]&H_in[909])^(data_in[142]&H_in[910])^(data_in[143]&H_in[911])^(data_in[144]&H_in[912])^(data_in[145]&H_in[913])^(data_in[146]&H_in[914])^(data_in[147]&H_in[915])^(data_in[148]&H_in[916])^(data_in[149]&H_in[917])^(data_in[150]&H_in[918])^(data_in[151]&H_in[919])^(data_in[152]&H_in[920])^(data_in[153]&H_in[921])^(data_in[154]&H_in[922])^(data_in[155]&H_in[923])^(data_in[156]&H_in[924])^(data_in[157]&H_in[925])^(data_in[158]&H_in[926])^(data_in[159]&H_in[927])^(data_in[160]&H_in[928])^(data_in[161]&H_in[929])^(data_in[162]&H_in[930])^(data_in[163]&H_in[931])^(data_in[164]&H_in[932])^(data_in[165]&H_in[933])^(data_in[166]&H_in[934])^(data_in[167]&H_in[935])^(data_in[168]&H_in[936])^(data_in[169]&H_in[937])^(data_in[170]&H_in[938])^(data_in[171]&H_in[939])^(data_in[172]&H_in[940])^(data_in[173]&H_in[941])^(data_in[174]&H_in[942])^(data_in[175]&H_in[943])^(data_in[176]&H_in[944])^(data_in[177]&H_in[945])^(data_in[178]&H_in[946])^(data_in[179]&H_in[947])^(data_in[180]&H_in[948])^(data_in[181]&H_in[949])^(data_in[182]&H_in[950])^(data_in[183]&H_in[951])^(data_in[184]&H_in[952])^(data_in[185]&H_in[953])^(data_in[186]&H_in[954])^(data_in[187]&H_in[955])^(data_in[188]&H_in[956])^(data_in[189]&H_in[957])^(data_in[190]&H_in[958])^(data_in[191]&H_in[959])^(data_in[192]&H_in[960])^(data_in[193]&H_in[961])^(data_in[194]&H_in[962])^(data_in[195]&H_in[963])^(data_in[196]&H_in[964])^(data_in[197]&H_in[965])^(data_in[198]&H_in[966])^(data_in[199]&H_in[967])^(data_in[200]&H_in[968])^(data_in[201]&H_in[969])^(data_in[202]&H_in[970])^(data_in[203]&H_in[971])^(data_in[204]&H_in[972])^(data_in[205]&H_in[973])^(data_in[206]&H_in[974])^(data_in[207]&H_in[975])^(data_in[208]&H_in[976])^(data_in[209]&H_in[977])^(data_in[210]&H_in[978])^(data_in[211]&H_in[979])^(data_in[212]&H_in[980])^(data_in[213]&H_in[981])^(data_in[214]&H_in[982])^(data_in[215]&H_in[983])^(data_in[216]&H_in[984])^(data_in[217]&H_in[985])^(data_in[218]&H_in[986])^(data_in[219]&H_in[987])^(data_in[220]&H_in[988])^(data_in[221]&H_in[989])^(data_in[222]&H_in[990])^(data_in[223]&H_in[991])^(data_in[224]&H_in[992])^(data_in[225]&H_in[993])^(data_in[226]&H_in[994])^(data_in[227]&H_in[995])^(data_in[228]&H_in[996])^(data_in[229]&H_in[997])^(data_in[230]&H_in[998])^(data_in[231]&H_in[999])^(data_in[232]&H_in[1000])^(data_in[233]&H_in[1001])^(data_in[234]&H_in[1002])^(data_in[235]&H_in[1003])^(data_in[236]&H_in[1004])^(data_in[237]&H_in[1005])^(data_in[238]&H_in[1006])^(data_in[239]&H_in[1007])^(data_in[240]&H_in[1008])^(data_in[241]&H_in[1009])^(data_in[242]&H_in[1010])^(data_in[243]&H_in[1011])^(data_in[244]&H_in[1012])^(data_in[245]&H_in[1013])^(data_in[246]&H_in[1014])^(data_in[247]&H_in[1015])^(data_in[248]&H_in[1016])^(data_in[249]&H_in[1017])^(data_in[250]&H_in[1018])^(data_in[251]&H_in[1019])^(data_in[252]&H_in[1020])^(data_in[253]&H_in[1021])^(data_in[254]&H_in[1022])^(data_in[255]&H_in[1023]);
         data_out[4]<=data_out[4]^(data_in[0]&H_in[1024])^(data_in[1]&H_in[1025])^(data_in[2]&H_in[1026])^(data_in[3]&H_in[1027])^(data_in[4]&H_in[1028])^(data_in[5]&H_in[1029])^(data_in[6]&H_in[1030])^(data_in[7]&H_in[1031])^(data_in[8]&H_in[1032])^(data_in[9]&H_in[1033])^(data_in[10]&H_in[1034])^(data_in[11]&H_in[1035])^(data_in[12]&H_in[1036])^(data_in[13]&H_in[1037])^(data_in[14]&H_in[1038])^(data_in[15]&H_in[1039])^(data_in[16]&H_in[1040])^(data_in[17]&H_in[1041])^(data_in[18]&H_in[1042])^(data_in[19]&H_in[1043])^(data_in[20]&H_in[1044])^(data_in[21]&H_in[1045])^(data_in[22]&H_in[1046])^(data_in[23]&H_in[1047])^(data_in[24]&H_in[1048])^(data_in[25]&H_in[1049])^(data_in[26]&H_in[1050])^(data_in[27]&H_in[1051])^(data_in[28]&H_in[1052])^(data_in[29]&H_in[1053])^(data_in[30]&H_in[1054])^(data_in[31]&H_in[1055])^(data_in[32]&H_in[1056])^(data_in[33]&H_in[1057])^(data_in[34]&H_in[1058])^(data_in[35]&H_in[1059])^(data_in[36]&H_in[1060])^(data_in[37]&H_in[1061])^(data_in[38]&H_in[1062])^(data_in[39]&H_in[1063])^(data_in[40]&H_in[1064])^(data_in[41]&H_in[1065])^(data_in[42]&H_in[1066])^(data_in[43]&H_in[1067])^(data_in[44]&H_in[1068])^(data_in[45]&H_in[1069])^(data_in[46]&H_in[1070])^(data_in[47]&H_in[1071])^(data_in[48]&H_in[1072])^(data_in[49]&H_in[1073])^(data_in[50]&H_in[1074])^(data_in[51]&H_in[1075])^(data_in[52]&H_in[1076])^(data_in[53]&H_in[1077])^(data_in[54]&H_in[1078])^(data_in[55]&H_in[1079])^(data_in[56]&H_in[1080])^(data_in[57]&H_in[1081])^(data_in[58]&H_in[1082])^(data_in[59]&H_in[1083])^(data_in[60]&H_in[1084])^(data_in[61]&H_in[1085])^(data_in[62]&H_in[1086])^(data_in[63]&H_in[1087])^(data_in[64]&H_in[1088])^(data_in[65]&H_in[1089])^(data_in[66]&H_in[1090])^(data_in[67]&H_in[1091])^(data_in[68]&H_in[1092])^(data_in[69]&H_in[1093])^(data_in[70]&H_in[1094])^(data_in[71]&H_in[1095])^(data_in[72]&H_in[1096])^(data_in[73]&H_in[1097])^(data_in[74]&H_in[1098])^(data_in[75]&H_in[1099])^(data_in[76]&H_in[1100])^(data_in[77]&H_in[1101])^(data_in[78]&H_in[1102])^(data_in[79]&H_in[1103])^(data_in[80]&H_in[1104])^(data_in[81]&H_in[1105])^(data_in[82]&H_in[1106])^(data_in[83]&H_in[1107])^(data_in[84]&H_in[1108])^(data_in[85]&H_in[1109])^(data_in[86]&H_in[1110])^(data_in[87]&H_in[1111])^(data_in[88]&H_in[1112])^(data_in[89]&H_in[1113])^(data_in[90]&H_in[1114])^(data_in[91]&H_in[1115])^(data_in[92]&H_in[1116])^(data_in[93]&H_in[1117])^(data_in[94]&H_in[1118])^(data_in[95]&H_in[1119])^(data_in[96]&H_in[1120])^(data_in[97]&H_in[1121])^(data_in[98]&H_in[1122])^(data_in[99]&H_in[1123])^(data_in[100]&H_in[1124])^(data_in[101]&H_in[1125])^(data_in[102]&H_in[1126])^(data_in[103]&H_in[1127])^(data_in[104]&H_in[1128])^(data_in[105]&H_in[1129])^(data_in[106]&H_in[1130])^(data_in[107]&H_in[1131])^(data_in[108]&H_in[1132])^(data_in[109]&H_in[1133])^(data_in[110]&H_in[1134])^(data_in[111]&H_in[1135])^(data_in[112]&H_in[1136])^(data_in[113]&H_in[1137])^(data_in[114]&H_in[1138])^(data_in[115]&H_in[1139])^(data_in[116]&H_in[1140])^(data_in[117]&H_in[1141])^(data_in[118]&H_in[1142])^(data_in[119]&H_in[1143])^(data_in[120]&H_in[1144])^(data_in[121]&H_in[1145])^(data_in[122]&H_in[1146])^(data_in[123]&H_in[1147])^(data_in[124]&H_in[1148])^(data_in[125]&H_in[1149])^(data_in[126]&H_in[1150])^(data_in[127]&H_in[1151])^(data_in[128]&H_in[1152])^(data_in[129]&H_in[1153])^(data_in[130]&H_in[1154])^(data_in[131]&H_in[1155])^(data_in[132]&H_in[1156])^(data_in[133]&H_in[1157])^(data_in[134]&H_in[1158])^(data_in[135]&H_in[1159])^(data_in[136]&H_in[1160])^(data_in[137]&H_in[1161])^(data_in[138]&H_in[1162])^(data_in[139]&H_in[1163])^(data_in[140]&H_in[1164])^(data_in[141]&H_in[1165])^(data_in[142]&H_in[1166])^(data_in[143]&H_in[1167])^(data_in[144]&H_in[1168])^(data_in[145]&H_in[1169])^(data_in[146]&H_in[1170])^(data_in[147]&H_in[1171])^(data_in[148]&H_in[1172])^(data_in[149]&H_in[1173])^(data_in[150]&H_in[1174])^(data_in[151]&H_in[1175])^(data_in[152]&H_in[1176])^(data_in[153]&H_in[1177])^(data_in[154]&H_in[1178])^(data_in[155]&H_in[1179])^(data_in[156]&H_in[1180])^(data_in[157]&H_in[1181])^(data_in[158]&H_in[1182])^(data_in[159]&H_in[1183])^(data_in[160]&H_in[1184])^(data_in[161]&H_in[1185])^(data_in[162]&H_in[1186])^(data_in[163]&H_in[1187])^(data_in[164]&H_in[1188])^(data_in[165]&H_in[1189])^(data_in[166]&H_in[1190])^(data_in[167]&H_in[1191])^(data_in[168]&H_in[1192])^(data_in[169]&H_in[1193])^(data_in[170]&H_in[1194])^(data_in[171]&H_in[1195])^(data_in[172]&H_in[1196])^(data_in[173]&H_in[1197])^(data_in[174]&H_in[1198])^(data_in[175]&H_in[1199])^(data_in[176]&H_in[1200])^(data_in[177]&H_in[1201])^(data_in[178]&H_in[1202])^(data_in[179]&H_in[1203])^(data_in[180]&H_in[1204])^(data_in[181]&H_in[1205])^(data_in[182]&H_in[1206])^(data_in[183]&H_in[1207])^(data_in[184]&H_in[1208])^(data_in[185]&H_in[1209])^(data_in[186]&H_in[1210])^(data_in[187]&H_in[1211])^(data_in[188]&H_in[1212])^(data_in[189]&H_in[1213])^(data_in[190]&H_in[1214])^(data_in[191]&H_in[1215])^(data_in[192]&H_in[1216])^(data_in[193]&H_in[1217])^(data_in[194]&H_in[1218])^(data_in[195]&H_in[1219])^(data_in[196]&H_in[1220])^(data_in[197]&H_in[1221])^(data_in[198]&H_in[1222])^(data_in[199]&H_in[1223])^(data_in[200]&H_in[1224])^(data_in[201]&H_in[1225])^(data_in[202]&H_in[1226])^(data_in[203]&H_in[1227])^(data_in[204]&H_in[1228])^(data_in[205]&H_in[1229])^(data_in[206]&H_in[1230])^(data_in[207]&H_in[1231])^(data_in[208]&H_in[1232])^(data_in[209]&H_in[1233])^(data_in[210]&H_in[1234])^(data_in[211]&H_in[1235])^(data_in[212]&H_in[1236])^(data_in[213]&H_in[1237])^(data_in[214]&H_in[1238])^(data_in[215]&H_in[1239])^(data_in[216]&H_in[1240])^(data_in[217]&H_in[1241])^(data_in[218]&H_in[1242])^(data_in[219]&H_in[1243])^(data_in[220]&H_in[1244])^(data_in[221]&H_in[1245])^(data_in[222]&H_in[1246])^(data_in[223]&H_in[1247])^(data_in[224]&H_in[1248])^(data_in[225]&H_in[1249])^(data_in[226]&H_in[1250])^(data_in[227]&H_in[1251])^(data_in[228]&H_in[1252])^(data_in[229]&H_in[1253])^(data_in[230]&H_in[1254])^(data_in[231]&H_in[1255])^(data_in[232]&H_in[1256])^(data_in[233]&H_in[1257])^(data_in[234]&H_in[1258])^(data_in[235]&H_in[1259])^(data_in[236]&H_in[1260])^(data_in[237]&H_in[1261])^(data_in[238]&H_in[1262])^(data_in[239]&H_in[1263])^(data_in[240]&H_in[1264])^(data_in[241]&H_in[1265])^(data_in[242]&H_in[1266])^(data_in[243]&H_in[1267])^(data_in[244]&H_in[1268])^(data_in[245]&H_in[1269])^(data_in[246]&H_in[1270])^(data_in[247]&H_in[1271])^(data_in[248]&H_in[1272])^(data_in[249]&H_in[1273])^(data_in[250]&H_in[1274])^(data_in[251]&H_in[1275])^(data_in[252]&H_in[1276])^(data_in[253]&H_in[1277])^(data_in[254]&H_in[1278])^(data_in[255]&H_in[1279]);
         data_out[5]<=data_out[5]^(data_in[0]&H_in[1280])^(data_in[1]&H_in[1281])^(data_in[2]&H_in[1282])^(data_in[3]&H_in[1283])^(data_in[4]&H_in[1284])^(data_in[5]&H_in[1285])^(data_in[6]&H_in[1286])^(data_in[7]&H_in[1287])^(data_in[8]&H_in[1288])^(data_in[9]&H_in[1289])^(data_in[10]&H_in[1290])^(data_in[11]&H_in[1291])^(data_in[12]&H_in[1292])^(data_in[13]&H_in[1293])^(data_in[14]&H_in[1294])^(data_in[15]&H_in[1295])^(data_in[16]&H_in[1296])^(data_in[17]&H_in[1297])^(data_in[18]&H_in[1298])^(data_in[19]&H_in[1299])^(data_in[20]&H_in[1300])^(data_in[21]&H_in[1301])^(data_in[22]&H_in[1302])^(data_in[23]&H_in[1303])^(data_in[24]&H_in[1304])^(data_in[25]&H_in[1305])^(data_in[26]&H_in[1306])^(data_in[27]&H_in[1307])^(data_in[28]&H_in[1308])^(data_in[29]&H_in[1309])^(data_in[30]&H_in[1310])^(data_in[31]&H_in[1311])^(data_in[32]&H_in[1312])^(data_in[33]&H_in[1313])^(data_in[34]&H_in[1314])^(data_in[35]&H_in[1315])^(data_in[36]&H_in[1316])^(data_in[37]&H_in[1317])^(data_in[38]&H_in[1318])^(data_in[39]&H_in[1319])^(data_in[40]&H_in[1320])^(data_in[41]&H_in[1321])^(data_in[42]&H_in[1322])^(data_in[43]&H_in[1323])^(data_in[44]&H_in[1324])^(data_in[45]&H_in[1325])^(data_in[46]&H_in[1326])^(data_in[47]&H_in[1327])^(data_in[48]&H_in[1328])^(data_in[49]&H_in[1329])^(data_in[50]&H_in[1330])^(data_in[51]&H_in[1331])^(data_in[52]&H_in[1332])^(data_in[53]&H_in[1333])^(data_in[54]&H_in[1334])^(data_in[55]&H_in[1335])^(data_in[56]&H_in[1336])^(data_in[57]&H_in[1337])^(data_in[58]&H_in[1338])^(data_in[59]&H_in[1339])^(data_in[60]&H_in[1340])^(data_in[61]&H_in[1341])^(data_in[62]&H_in[1342])^(data_in[63]&H_in[1343])^(data_in[64]&H_in[1344])^(data_in[65]&H_in[1345])^(data_in[66]&H_in[1346])^(data_in[67]&H_in[1347])^(data_in[68]&H_in[1348])^(data_in[69]&H_in[1349])^(data_in[70]&H_in[1350])^(data_in[71]&H_in[1351])^(data_in[72]&H_in[1352])^(data_in[73]&H_in[1353])^(data_in[74]&H_in[1354])^(data_in[75]&H_in[1355])^(data_in[76]&H_in[1356])^(data_in[77]&H_in[1357])^(data_in[78]&H_in[1358])^(data_in[79]&H_in[1359])^(data_in[80]&H_in[1360])^(data_in[81]&H_in[1361])^(data_in[82]&H_in[1362])^(data_in[83]&H_in[1363])^(data_in[84]&H_in[1364])^(data_in[85]&H_in[1365])^(data_in[86]&H_in[1366])^(data_in[87]&H_in[1367])^(data_in[88]&H_in[1368])^(data_in[89]&H_in[1369])^(data_in[90]&H_in[1370])^(data_in[91]&H_in[1371])^(data_in[92]&H_in[1372])^(data_in[93]&H_in[1373])^(data_in[94]&H_in[1374])^(data_in[95]&H_in[1375])^(data_in[96]&H_in[1376])^(data_in[97]&H_in[1377])^(data_in[98]&H_in[1378])^(data_in[99]&H_in[1379])^(data_in[100]&H_in[1380])^(data_in[101]&H_in[1381])^(data_in[102]&H_in[1382])^(data_in[103]&H_in[1383])^(data_in[104]&H_in[1384])^(data_in[105]&H_in[1385])^(data_in[106]&H_in[1386])^(data_in[107]&H_in[1387])^(data_in[108]&H_in[1388])^(data_in[109]&H_in[1389])^(data_in[110]&H_in[1390])^(data_in[111]&H_in[1391])^(data_in[112]&H_in[1392])^(data_in[113]&H_in[1393])^(data_in[114]&H_in[1394])^(data_in[115]&H_in[1395])^(data_in[116]&H_in[1396])^(data_in[117]&H_in[1397])^(data_in[118]&H_in[1398])^(data_in[119]&H_in[1399])^(data_in[120]&H_in[1400])^(data_in[121]&H_in[1401])^(data_in[122]&H_in[1402])^(data_in[123]&H_in[1403])^(data_in[124]&H_in[1404])^(data_in[125]&H_in[1405])^(data_in[126]&H_in[1406])^(data_in[127]&H_in[1407])^(data_in[128]&H_in[1408])^(data_in[129]&H_in[1409])^(data_in[130]&H_in[1410])^(data_in[131]&H_in[1411])^(data_in[132]&H_in[1412])^(data_in[133]&H_in[1413])^(data_in[134]&H_in[1414])^(data_in[135]&H_in[1415])^(data_in[136]&H_in[1416])^(data_in[137]&H_in[1417])^(data_in[138]&H_in[1418])^(data_in[139]&H_in[1419])^(data_in[140]&H_in[1420])^(data_in[141]&H_in[1421])^(data_in[142]&H_in[1422])^(data_in[143]&H_in[1423])^(data_in[144]&H_in[1424])^(data_in[145]&H_in[1425])^(data_in[146]&H_in[1426])^(data_in[147]&H_in[1427])^(data_in[148]&H_in[1428])^(data_in[149]&H_in[1429])^(data_in[150]&H_in[1430])^(data_in[151]&H_in[1431])^(data_in[152]&H_in[1432])^(data_in[153]&H_in[1433])^(data_in[154]&H_in[1434])^(data_in[155]&H_in[1435])^(data_in[156]&H_in[1436])^(data_in[157]&H_in[1437])^(data_in[158]&H_in[1438])^(data_in[159]&H_in[1439])^(data_in[160]&H_in[1440])^(data_in[161]&H_in[1441])^(data_in[162]&H_in[1442])^(data_in[163]&H_in[1443])^(data_in[164]&H_in[1444])^(data_in[165]&H_in[1445])^(data_in[166]&H_in[1446])^(data_in[167]&H_in[1447])^(data_in[168]&H_in[1448])^(data_in[169]&H_in[1449])^(data_in[170]&H_in[1450])^(data_in[171]&H_in[1451])^(data_in[172]&H_in[1452])^(data_in[173]&H_in[1453])^(data_in[174]&H_in[1454])^(data_in[175]&H_in[1455])^(data_in[176]&H_in[1456])^(data_in[177]&H_in[1457])^(data_in[178]&H_in[1458])^(data_in[179]&H_in[1459])^(data_in[180]&H_in[1460])^(data_in[181]&H_in[1461])^(data_in[182]&H_in[1462])^(data_in[183]&H_in[1463])^(data_in[184]&H_in[1464])^(data_in[185]&H_in[1465])^(data_in[186]&H_in[1466])^(data_in[187]&H_in[1467])^(data_in[188]&H_in[1468])^(data_in[189]&H_in[1469])^(data_in[190]&H_in[1470])^(data_in[191]&H_in[1471])^(data_in[192]&H_in[1472])^(data_in[193]&H_in[1473])^(data_in[194]&H_in[1474])^(data_in[195]&H_in[1475])^(data_in[196]&H_in[1476])^(data_in[197]&H_in[1477])^(data_in[198]&H_in[1478])^(data_in[199]&H_in[1479])^(data_in[200]&H_in[1480])^(data_in[201]&H_in[1481])^(data_in[202]&H_in[1482])^(data_in[203]&H_in[1483])^(data_in[204]&H_in[1484])^(data_in[205]&H_in[1485])^(data_in[206]&H_in[1486])^(data_in[207]&H_in[1487])^(data_in[208]&H_in[1488])^(data_in[209]&H_in[1489])^(data_in[210]&H_in[1490])^(data_in[211]&H_in[1491])^(data_in[212]&H_in[1492])^(data_in[213]&H_in[1493])^(data_in[214]&H_in[1494])^(data_in[215]&H_in[1495])^(data_in[216]&H_in[1496])^(data_in[217]&H_in[1497])^(data_in[218]&H_in[1498])^(data_in[219]&H_in[1499])^(data_in[220]&H_in[1500])^(data_in[221]&H_in[1501])^(data_in[222]&H_in[1502])^(data_in[223]&H_in[1503])^(data_in[224]&H_in[1504])^(data_in[225]&H_in[1505])^(data_in[226]&H_in[1506])^(data_in[227]&H_in[1507])^(data_in[228]&H_in[1508])^(data_in[229]&H_in[1509])^(data_in[230]&H_in[1510])^(data_in[231]&H_in[1511])^(data_in[232]&H_in[1512])^(data_in[233]&H_in[1513])^(data_in[234]&H_in[1514])^(data_in[235]&H_in[1515])^(data_in[236]&H_in[1516])^(data_in[237]&H_in[1517])^(data_in[238]&H_in[1518])^(data_in[239]&H_in[1519])^(data_in[240]&H_in[1520])^(data_in[241]&H_in[1521])^(data_in[242]&H_in[1522])^(data_in[243]&H_in[1523])^(data_in[244]&H_in[1524])^(data_in[245]&H_in[1525])^(data_in[246]&H_in[1526])^(data_in[247]&H_in[1527])^(data_in[248]&H_in[1528])^(data_in[249]&H_in[1529])^(data_in[250]&H_in[1530])^(data_in[251]&H_in[1531])^(data_in[252]&H_in[1532])^(data_in[253]&H_in[1533])^(data_in[254]&H_in[1534])^(data_in[255]&H_in[1535]);
         data_out[6]<=data_out[6]^(data_in[0]&H_in[1536])^(data_in[1]&H_in[1537])^(data_in[2]&H_in[1538])^(data_in[3]&H_in[1539])^(data_in[4]&H_in[1540])^(data_in[5]&H_in[1541])^(data_in[6]&H_in[1542])^(data_in[7]&H_in[1543])^(data_in[8]&H_in[1544])^(data_in[9]&H_in[1545])^(data_in[10]&H_in[1546])^(data_in[11]&H_in[1547])^(data_in[12]&H_in[1548])^(data_in[13]&H_in[1549])^(data_in[14]&H_in[1550])^(data_in[15]&H_in[1551])^(data_in[16]&H_in[1552])^(data_in[17]&H_in[1553])^(data_in[18]&H_in[1554])^(data_in[19]&H_in[1555])^(data_in[20]&H_in[1556])^(data_in[21]&H_in[1557])^(data_in[22]&H_in[1558])^(data_in[23]&H_in[1559])^(data_in[24]&H_in[1560])^(data_in[25]&H_in[1561])^(data_in[26]&H_in[1562])^(data_in[27]&H_in[1563])^(data_in[28]&H_in[1564])^(data_in[29]&H_in[1565])^(data_in[30]&H_in[1566])^(data_in[31]&H_in[1567])^(data_in[32]&H_in[1568])^(data_in[33]&H_in[1569])^(data_in[34]&H_in[1570])^(data_in[35]&H_in[1571])^(data_in[36]&H_in[1572])^(data_in[37]&H_in[1573])^(data_in[38]&H_in[1574])^(data_in[39]&H_in[1575])^(data_in[40]&H_in[1576])^(data_in[41]&H_in[1577])^(data_in[42]&H_in[1578])^(data_in[43]&H_in[1579])^(data_in[44]&H_in[1580])^(data_in[45]&H_in[1581])^(data_in[46]&H_in[1582])^(data_in[47]&H_in[1583])^(data_in[48]&H_in[1584])^(data_in[49]&H_in[1585])^(data_in[50]&H_in[1586])^(data_in[51]&H_in[1587])^(data_in[52]&H_in[1588])^(data_in[53]&H_in[1589])^(data_in[54]&H_in[1590])^(data_in[55]&H_in[1591])^(data_in[56]&H_in[1592])^(data_in[57]&H_in[1593])^(data_in[58]&H_in[1594])^(data_in[59]&H_in[1595])^(data_in[60]&H_in[1596])^(data_in[61]&H_in[1597])^(data_in[62]&H_in[1598])^(data_in[63]&H_in[1599])^(data_in[64]&H_in[1600])^(data_in[65]&H_in[1601])^(data_in[66]&H_in[1602])^(data_in[67]&H_in[1603])^(data_in[68]&H_in[1604])^(data_in[69]&H_in[1605])^(data_in[70]&H_in[1606])^(data_in[71]&H_in[1607])^(data_in[72]&H_in[1608])^(data_in[73]&H_in[1609])^(data_in[74]&H_in[1610])^(data_in[75]&H_in[1611])^(data_in[76]&H_in[1612])^(data_in[77]&H_in[1613])^(data_in[78]&H_in[1614])^(data_in[79]&H_in[1615])^(data_in[80]&H_in[1616])^(data_in[81]&H_in[1617])^(data_in[82]&H_in[1618])^(data_in[83]&H_in[1619])^(data_in[84]&H_in[1620])^(data_in[85]&H_in[1621])^(data_in[86]&H_in[1622])^(data_in[87]&H_in[1623])^(data_in[88]&H_in[1624])^(data_in[89]&H_in[1625])^(data_in[90]&H_in[1626])^(data_in[91]&H_in[1627])^(data_in[92]&H_in[1628])^(data_in[93]&H_in[1629])^(data_in[94]&H_in[1630])^(data_in[95]&H_in[1631])^(data_in[96]&H_in[1632])^(data_in[97]&H_in[1633])^(data_in[98]&H_in[1634])^(data_in[99]&H_in[1635])^(data_in[100]&H_in[1636])^(data_in[101]&H_in[1637])^(data_in[102]&H_in[1638])^(data_in[103]&H_in[1639])^(data_in[104]&H_in[1640])^(data_in[105]&H_in[1641])^(data_in[106]&H_in[1642])^(data_in[107]&H_in[1643])^(data_in[108]&H_in[1644])^(data_in[109]&H_in[1645])^(data_in[110]&H_in[1646])^(data_in[111]&H_in[1647])^(data_in[112]&H_in[1648])^(data_in[113]&H_in[1649])^(data_in[114]&H_in[1650])^(data_in[115]&H_in[1651])^(data_in[116]&H_in[1652])^(data_in[117]&H_in[1653])^(data_in[118]&H_in[1654])^(data_in[119]&H_in[1655])^(data_in[120]&H_in[1656])^(data_in[121]&H_in[1657])^(data_in[122]&H_in[1658])^(data_in[123]&H_in[1659])^(data_in[124]&H_in[1660])^(data_in[125]&H_in[1661])^(data_in[126]&H_in[1662])^(data_in[127]&H_in[1663])^(data_in[128]&H_in[1664])^(data_in[129]&H_in[1665])^(data_in[130]&H_in[1666])^(data_in[131]&H_in[1667])^(data_in[132]&H_in[1668])^(data_in[133]&H_in[1669])^(data_in[134]&H_in[1670])^(data_in[135]&H_in[1671])^(data_in[136]&H_in[1672])^(data_in[137]&H_in[1673])^(data_in[138]&H_in[1674])^(data_in[139]&H_in[1675])^(data_in[140]&H_in[1676])^(data_in[141]&H_in[1677])^(data_in[142]&H_in[1678])^(data_in[143]&H_in[1679])^(data_in[144]&H_in[1680])^(data_in[145]&H_in[1681])^(data_in[146]&H_in[1682])^(data_in[147]&H_in[1683])^(data_in[148]&H_in[1684])^(data_in[149]&H_in[1685])^(data_in[150]&H_in[1686])^(data_in[151]&H_in[1687])^(data_in[152]&H_in[1688])^(data_in[153]&H_in[1689])^(data_in[154]&H_in[1690])^(data_in[155]&H_in[1691])^(data_in[156]&H_in[1692])^(data_in[157]&H_in[1693])^(data_in[158]&H_in[1694])^(data_in[159]&H_in[1695])^(data_in[160]&H_in[1696])^(data_in[161]&H_in[1697])^(data_in[162]&H_in[1698])^(data_in[163]&H_in[1699])^(data_in[164]&H_in[1700])^(data_in[165]&H_in[1701])^(data_in[166]&H_in[1702])^(data_in[167]&H_in[1703])^(data_in[168]&H_in[1704])^(data_in[169]&H_in[1705])^(data_in[170]&H_in[1706])^(data_in[171]&H_in[1707])^(data_in[172]&H_in[1708])^(data_in[173]&H_in[1709])^(data_in[174]&H_in[1710])^(data_in[175]&H_in[1711])^(data_in[176]&H_in[1712])^(data_in[177]&H_in[1713])^(data_in[178]&H_in[1714])^(data_in[179]&H_in[1715])^(data_in[180]&H_in[1716])^(data_in[181]&H_in[1717])^(data_in[182]&H_in[1718])^(data_in[183]&H_in[1719])^(data_in[184]&H_in[1720])^(data_in[185]&H_in[1721])^(data_in[186]&H_in[1722])^(data_in[187]&H_in[1723])^(data_in[188]&H_in[1724])^(data_in[189]&H_in[1725])^(data_in[190]&H_in[1726])^(data_in[191]&H_in[1727])^(data_in[192]&H_in[1728])^(data_in[193]&H_in[1729])^(data_in[194]&H_in[1730])^(data_in[195]&H_in[1731])^(data_in[196]&H_in[1732])^(data_in[197]&H_in[1733])^(data_in[198]&H_in[1734])^(data_in[199]&H_in[1735])^(data_in[200]&H_in[1736])^(data_in[201]&H_in[1737])^(data_in[202]&H_in[1738])^(data_in[203]&H_in[1739])^(data_in[204]&H_in[1740])^(data_in[205]&H_in[1741])^(data_in[206]&H_in[1742])^(data_in[207]&H_in[1743])^(data_in[208]&H_in[1744])^(data_in[209]&H_in[1745])^(data_in[210]&H_in[1746])^(data_in[211]&H_in[1747])^(data_in[212]&H_in[1748])^(data_in[213]&H_in[1749])^(data_in[214]&H_in[1750])^(data_in[215]&H_in[1751])^(data_in[216]&H_in[1752])^(data_in[217]&H_in[1753])^(data_in[218]&H_in[1754])^(data_in[219]&H_in[1755])^(data_in[220]&H_in[1756])^(data_in[221]&H_in[1757])^(data_in[222]&H_in[1758])^(data_in[223]&H_in[1759])^(data_in[224]&H_in[1760])^(data_in[225]&H_in[1761])^(data_in[226]&H_in[1762])^(data_in[227]&H_in[1763])^(data_in[228]&H_in[1764])^(data_in[229]&H_in[1765])^(data_in[230]&H_in[1766])^(data_in[231]&H_in[1767])^(data_in[232]&H_in[1768])^(data_in[233]&H_in[1769])^(data_in[234]&H_in[1770])^(data_in[235]&H_in[1771])^(data_in[236]&H_in[1772])^(data_in[237]&H_in[1773])^(data_in[238]&H_in[1774])^(data_in[239]&H_in[1775])^(data_in[240]&H_in[1776])^(data_in[241]&H_in[1777])^(data_in[242]&H_in[1778])^(data_in[243]&H_in[1779])^(data_in[244]&H_in[1780])^(data_in[245]&H_in[1781])^(data_in[246]&H_in[1782])^(data_in[247]&H_in[1783])^(data_in[248]&H_in[1784])^(data_in[249]&H_in[1785])^(data_in[250]&H_in[1786])^(data_in[251]&H_in[1787])^(data_in[252]&H_in[1788])^(data_in[253]&H_in[1789])^(data_in[254]&H_in[1790])^(data_in[255]&H_in[1791]);
         data_out[7]<=data_out[7]^(data_in[0]&H_in[1792])^(data_in[1]&H_in[1793])^(data_in[2]&H_in[1794])^(data_in[3]&H_in[1795])^(data_in[4]&H_in[1796])^(data_in[5]&H_in[1797])^(data_in[6]&H_in[1798])^(data_in[7]&H_in[1799])^(data_in[8]&H_in[1800])^(data_in[9]&H_in[1801])^(data_in[10]&H_in[1802])^(data_in[11]&H_in[1803])^(data_in[12]&H_in[1804])^(data_in[13]&H_in[1805])^(data_in[14]&H_in[1806])^(data_in[15]&H_in[1807])^(data_in[16]&H_in[1808])^(data_in[17]&H_in[1809])^(data_in[18]&H_in[1810])^(data_in[19]&H_in[1811])^(data_in[20]&H_in[1812])^(data_in[21]&H_in[1813])^(data_in[22]&H_in[1814])^(data_in[23]&H_in[1815])^(data_in[24]&H_in[1816])^(data_in[25]&H_in[1817])^(data_in[26]&H_in[1818])^(data_in[27]&H_in[1819])^(data_in[28]&H_in[1820])^(data_in[29]&H_in[1821])^(data_in[30]&H_in[1822])^(data_in[31]&H_in[1823])^(data_in[32]&H_in[1824])^(data_in[33]&H_in[1825])^(data_in[34]&H_in[1826])^(data_in[35]&H_in[1827])^(data_in[36]&H_in[1828])^(data_in[37]&H_in[1829])^(data_in[38]&H_in[1830])^(data_in[39]&H_in[1831])^(data_in[40]&H_in[1832])^(data_in[41]&H_in[1833])^(data_in[42]&H_in[1834])^(data_in[43]&H_in[1835])^(data_in[44]&H_in[1836])^(data_in[45]&H_in[1837])^(data_in[46]&H_in[1838])^(data_in[47]&H_in[1839])^(data_in[48]&H_in[1840])^(data_in[49]&H_in[1841])^(data_in[50]&H_in[1842])^(data_in[51]&H_in[1843])^(data_in[52]&H_in[1844])^(data_in[53]&H_in[1845])^(data_in[54]&H_in[1846])^(data_in[55]&H_in[1847])^(data_in[56]&H_in[1848])^(data_in[57]&H_in[1849])^(data_in[58]&H_in[1850])^(data_in[59]&H_in[1851])^(data_in[60]&H_in[1852])^(data_in[61]&H_in[1853])^(data_in[62]&H_in[1854])^(data_in[63]&H_in[1855])^(data_in[64]&H_in[1856])^(data_in[65]&H_in[1857])^(data_in[66]&H_in[1858])^(data_in[67]&H_in[1859])^(data_in[68]&H_in[1860])^(data_in[69]&H_in[1861])^(data_in[70]&H_in[1862])^(data_in[71]&H_in[1863])^(data_in[72]&H_in[1864])^(data_in[73]&H_in[1865])^(data_in[74]&H_in[1866])^(data_in[75]&H_in[1867])^(data_in[76]&H_in[1868])^(data_in[77]&H_in[1869])^(data_in[78]&H_in[1870])^(data_in[79]&H_in[1871])^(data_in[80]&H_in[1872])^(data_in[81]&H_in[1873])^(data_in[82]&H_in[1874])^(data_in[83]&H_in[1875])^(data_in[84]&H_in[1876])^(data_in[85]&H_in[1877])^(data_in[86]&H_in[1878])^(data_in[87]&H_in[1879])^(data_in[88]&H_in[1880])^(data_in[89]&H_in[1881])^(data_in[90]&H_in[1882])^(data_in[91]&H_in[1883])^(data_in[92]&H_in[1884])^(data_in[93]&H_in[1885])^(data_in[94]&H_in[1886])^(data_in[95]&H_in[1887])^(data_in[96]&H_in[1888])^(data_in[97]&H_in[1889])^(data_in[98]&H_in[1890])^(data_in[99]&H_in[1891])^(data_in[100]&H_in[1892])^(data_in[101]&H_in[1893])^(data_in[102]&H_in[1894])^(data_in[103]&H_in[1895])^(data_in[104]&H_in[1896])^(data_in[105]&H_in[1897])^(data_in[106]&H_in[1898])^(data_in[107]&H_in[1899])^(data_in[108]&H_in[1900])^(data_in[109]&H_in[1901])^(data_in[110]&H_in[1902])^(data_in[111]&H_in[1903])^(data_in[112]&H_in[1904])^(data_in[113]&H_in[1905])^(data_in[114]&H_in[1906])^(data_in[115]&H_in[1907])^(data_in[116]&H_in[1908])^(data_in[117]&H_in[1909])^(data_in[118]&H_in[1910])^(data_in[119]&H_in[1911])^(data_in[120]&H_in[1912])^(data_in[121]&H_in[1913])^(data_in[122]&H_in[1914])^(data_in[123]&H_in[1915])^(data_in[124]&H_in[1916])^(data_in[125]&H_in[1917])^(data_in[126]&H_in[1918])^(data_in[127]&H_in[1919])^(data_in[128]&H_in[1920])^(data_in[129]&H_in[1921])^(data_in[130]&H_in[1922])^(data_in[131]&H_in[1923])^(data_in[132]&H_in[1924])^(data_in[133]&H_in[1925])^(data_in[134]&H_in[1926])^(data_in[135]&H_in[1927])^(data_in[136]&H_in[1928])^(data_in[137]&H_in[1929])^(data_in[138]&H_in[1930])^(data_in[139]&H_in[1931])^(data_in[140]&H_in[1932])^(data_in[141]&H_in[1933])^(data_in[142]&H_in[1934])^(data_in[143]&H_in[1935])^(data_in[144]&H_in[1936])^(data_in[145]&H_in[1937])^(data_in[146]&H_in[1938])^(data_in[147]&H_in[1939])^(data_in[148]&H_in[1940])^(data_in[149]&H_in[1941])^(data_in[150]&H_in[1942])^(data_in[151]&H_in[1943])^(data_in[152]&H_in[1944])^(data_in[153]&H_in[1945])^(data_in[154]&H_in[1946])^(data_in[155]&H_in[1947])^(data_in[156]&H_in[1948])^(data_in[157]&H_in[1949])^(data_in[158]&H_in[1950])^(data_in[159]&H_in[1951])^(data_in[160]&H_in[1952])^(data_in[161]&H_in[1953])^(data_in[162]&H_in[1954])^(data_in[163]&H_in[1955])^(data_in[164]&H_in[1956])^(data_in[165]&H_in[1957])^(data_in[166]&H_in[1958])^(data_in[167]&H_in[1959])^(data_in[168]&H_in[1960])^(data_in[169]&H_in[1961])^(data_in[170]&H_in[1962])^(data_in[171]&H_in[1963])^(data_in[172]&H_in[1964])^(data_in[173]&H_in[1965])^(data_in[174]&H_in[1966])^(data_in[175]&H_in[1967])^(data_in[176]&H_in[1968])^(data_in[177]&H_in[1969])^(data_in[178]&H_in[1970])^(data_in[179]&H_in[1971])^(data_in[180]&H_in[1972])^(data_in[181]&H_in[1973])^(data_in[182]&H_in[1974])^(data_in[183]&H_in[1975])^(data_in[184]&H_in[1976])^(data_in[185]&H_in[1977])^(data_in[186]&H_in[1978])^(data_in[187]&H_in[1979])^(data_in[188]&H_in[1980])^(data_in[189]&H_in[1981])^(data_in[190]&H_in[1982])^(data_in[191]&H_in[1983])^(data_in[192]&H_in[1984])^(data_in[193]&H_in[1985])^(data_in[194]&H_in[1986])^(data_in[195]&H_in[1987])^(data_in[196]&H_in[1988])^(data_in[197]&H_in[1989])^(data_in[198]&H_in[1990])^(data_in[199]&H_in[1991])^(data_in[200]&H_in[1992])^(data_in[201]&H_in[1993])^(data_in[202]&H_in[1994])^(data_in[203]&H_in[1995])^(data_in[204]&H_in[1996])^(data_in[205]&H_in[1997])^(data_in[206]&H_in[1998])^(data_in[207]&H_in[1999])^(data_in[208]&H_in[2000])^(data_in[209]&H_in[2001])^(data_in[210]&H_in[2002])^(data_in[211]&H_in[2003])^(data_in[212]&H_in[2004])^(data_in[213]&H_in[2005])^(data_in[214]&H_in[2006])^(data_in[215]&H_in[2007])^(data_in[216]&H_in[2008])^(data_in[217]&H_in[2009])^(data_in[218]&H_in[2010])^(data_in[219]&H_in[2011])^(data_in[220]&H_in[2012])^(data_in[221]&H_in[2013])^(data_in[222]&H_in[2014])^(data_in[223]&H_in[2015])^(data_in[224]&H_in[2016])^(data_in[225]&H_in[2017])^(data_in[226]&H_in[2018])^(data_in[227]&H_in[2019])^(data_in[228]&H_in[2020])^(data_in[229]&H_in[2021])^(data_in[230]&H_in[2022])^(data_in[231]&H_in[2023])^(data_in[232]&H_in[2024])^(data_in[233]&H_in[2025])^(data_in[234]&H_in[2026])^(data_in[235]&H_in[2027])^(data_in[236]&H_in[2028])^(data_in[237]&H_in[2029])^(data_in[238]&H_in[2030])^(data_in[239]&H_in[2031])^(data_in[240]&H_in[2032])^(data_in[241]&H_in[2033])^(data_in[242]&H_in[2034])^(data_in[243]&H_in[2035])^(data_in[244]&H_in[2036])^(data_in[245]&H_in[2037])^(data_in[246]&H_in[2038])^(data_in[247]&H_in[2039])^(data_in[248]&H_in[2040])^(data_in[249]&H_in[2041])^(data_in[250]&H_in[2042])^(data_in[251]&H_in[2043])^(data_in[252]&H_in[2044])^(data_in[253]&H_in[2045])^(data_in[254]&H_in[2046])^(data_in[255]&H_in[2047]);
         data_out[8]<=data_out[8]^(data_in[0]&H_in[2048])^(data_in[1]&H_in[2049])^(data_in[2]&H_in[2050])^(data_in[3]&H_in[2051])^(data_in[4]&H_in[2052])^(data_in[5]&H_in[2053])^(data_in[6]&H_in[2054])^(data_in[7]&H_in[2055])^(data_in[8]&H_in[2056])^(data_in[9]&H_in[2057])^(data_in[10]&H_in[2058])^(data_in[11]&H_in[2059])^(data_in[12]&H_in[2060])^(data_in[13]&H_in[2061])^(data_in[14]&H_in[2062])^(data_in[15]&H_in[2063])^(data_in[16]&H_in[2064])^(data_in[17]&H_in[2065])^(data_in[18]&H_in[2066])^(data_in[19]&H_in[2067])^(data_in[20]&H_in[2068])^(data_in[21]&H_in[2069])^(data_in[22]&H_in[2070])^(data_in[23]&H_in[2071])^(data_in[24]&H_in[2072])^(data_in[25]&H_in[2073])^(data_in[26]&H_in[2074])^(data_in[27]&H_in[2075])^(data_in[28]&H_in[2076])^(data_in[29]&H_in[2077])^(data_in[30]&H_in[2078])^(data_in[31]&H_in[2079])^(data_in[32]&H_in[2080])^(data_in[33]&H_in[2081])^(data_in[34]&H_in[2082])^(data_in[35]&H_in[2083])^(data_in[36]&H_in[2084])^(data_in[37]&H_in[2085])^(data_in[38]&H_in[2086])^(data_in[39]&H_in[2087])^(data_in[40]&H_in[2088])^(data_in[41]&H_in[2089])^(data_in[42]&H_in[2090])^(data_in[43]&H_in[2091])^(data_in[44]&H_in[2092])^(data_in[45]&H_in[2093])^(data_in[46]&H_in[2094])^(data_in[47]&H_in[2095])^(data_in[48]&H_in[2096])^(data_in[49]&H_in[2097])^(data_in[50]&H_in[2098])^(data_in[51]&H_in[2099])^(data_in[52]&H_in[2100])^(data_in[53]&H_in[2101])^(data_in[54]&H_in[2102])^(data_in[55]&H_in[2103])^(data_in[56]&H_in[2104])^(data_in[57]&H_in[2105])^(data_in[58]&H_in[2106])^(data_in[59]&H_in[2107])^(data_in[60]&H_in[2108])^(data_in[61]&H_in[2109])^(data_in[62]&H_in[2110])^(data_in[63]&H_in[2111])^(data_in[64]&H_in[2112])^(data_in[65]&H_in[2113])^(data_in[66]&H_in[2114])^(data_in[67]&H_in[2115])^(data_in[68]&H_in[2116])^(data_in[69]&H_in[2117])^(data_in[70]&H_in[2118])^(data_in[71]&H_in[2119])^(data_in[72]&H_in[2120])^(data_in[73]&H_in[2121])^(data_in[74]&H_in[2122])^(data_in[75]&H_in[2123])^(data_in[76]&H_in[2124])^(data_in[77]&H_in[2125])^(data_in[78]&H_in[2126])^(data_in[79]&H_in[2127])^(data_in[80]&H_in[2128])^(data_in[81]&H_in[2129])^(data_in[82]&H_in[2130])^(data_in[83]&H_in[2131])^(data_in[84]&H_in[2132])^(data_in[85]&H_in[2133])^(data_in[86]&H_in[2134])^(data_in[87]&H_in[2135])^(data_in[88]&H_in[2136])^(data_in[89]&H_in[2137])^(data_in[90]&H_in[2138])^(data_in[91]&H_in[2139])^(data_in[92]&H_in[2140])^(data_in[93]&H_in[2141])^(data_in[94]&H_in[2142])^(data_in[95]&H_in[2143])^(data_in[96]&H_in[2144])^(data_in[97]&H_in[2145])^(data_in[98]&H_in[2146])^(data_in[99]&H_in[2147])^(data_in[100]&H_in[2148])^(data_in[101]&H_in[2149])^(data_in[102]&H_in[2150])^(data_in[103]&H_in[2151])^(data_in[104]&H_in[2152])^(data_in[105]&H_in[2153])^(data_in[106]&H_in[2154])^(data_in[107]&H_in[2155])^(data_in[108]&H_in[2156])^(data_in[109]&H_in[2157])^(data_in[110]&H_in[2158])^(data_in[111]&H_in[2159])^(data_in[112]&H_in[2160])^(data_in[113]&H_in[2161])^(data_in[114]&H_in[2162])^(data_in[115]&H_in[2163])^(data_in[116]&H_in[2164])^(data_in[117]&H_in[2165])^(data_in[118]&H_in[2166])^(data_in[119]&H_in[2167])^(data_in[120]&H_in[2168])^(data_in[121]&H_in[2169])^(data_in[122]&H_in[2170])^(data_in[123]&H_in[2171])^(data_in[124]&H_in[2172])^(data_in[125]&H_in[2173])^(data_in[126]&H_in[2174])^(data_in[127]&H_in[2175])^(data_in[128]&H_in[2176])^(data_in[129]&H_in[2177])^(data_in[130]&H_in[2178])^(data_in[131]&H_in[2179])^(data_in[132]&H_in[2180])^(data_in[133]&H_in[2181])^(data_in[134]&H_in[2182])^(data_in[135]&H_in[2183])^(data_in[136]&H_in[2184])^(data_in[137]&H_in[2185])^(data_in[138]&H_in[2186])^(data_in[139]&H_in[2187])^(data_in[140]&H_in[2188])^(data_in[141]&H_in[2189])^(data_in[142]&H_in[2190])^(data_in[143]&H_in[2191])^(data_in[144]&H_in[2192])^(data_in[145]&H_in[2193])^(data_in[146]&H_in[2194])^(data_in[147]&H_in[2195])^(data_in[148]&H_in[2196])^(data_in[149]&H_in[2197])^(data_in[150]&H_in[2198])^(data_in[151]&H_in[2199])^(data_in[152]&H_in[2200])^(data_in[153]&H_in[2201])^(data_in[154]&H_in[2202])^(data_in[155]&H_in[2203])^(data_in[156]&H_in[2204])^(data_in[157]&H_in[2205])^(data_in[158]&H_in[2206])^(data_in[159]&H_in[2207])^(data_in[160]&H_in[2208])^(data_in[161]&H_in[2209])^(data_in[162]&H_in[2210])^(data_in[163]&H_in[2211])^(data_in[164]&H_in[2212])^(data_in[165]&H_in[2213])^(data_in[166]&H_in[2214])^(data_in[167]&H_in[2215])^(data_in[168]&H_in[2216])^(data_in[169]&H_in[2217])^(data_in[170]&H_in[2218])^(data_in[171]&H_in[2219])^(data_in[172]&H_in[2220])^(data_in[173]&H_in[2221])^(data_in[174]&H_in[2222])^(data_in[175]&H_in[2223])^(data_in[176]&H_in[2224])^(data_in[177]&H_in[2225])^(data_in[178]&H_in[2226])^(data_in[179]&H_in[2227])^(data_in[180]&H_in[2228])^(data_in[181]&H_in[2229])^(data_in[182]&H_in[2230])^(data_in[183]&H_in[2231])^(data_in[184]&H_in[2232])^(data_in[185]&H_in[2233])^(data_in[186]&H_in[2234])^(data_in[187]&H_in[2235])^(data_in[188]&H_in[2236])^(data_in[189]&H_in[2237])^(data_in[190]&H_in[2238])^(data_in[191]&H_in[2239])^(data_in[192]&H_in[2240])^(data_in[193]&H_in[2241])^(data_in[194]&H_in[2242])^(data_in[195]&H_in[2243])^(data_in[196]&H_in[2244])^(data_in[197]&H_in[2245])^(data_in[198]&H_in[2246])^(data_in[199]&H_in[2247])^(data_in[200]&H_in[2248])^(data_in[201]&H_in[2249])^(data_in[202]&H_in[2250])^(data_in[203]&H_in[2251])^(data_in[204]&H_in[2252])^(data_in[205]&H_in[2253])^(data_in[206]&H_in[2254])^(data_in[207]&H_in[2255])^(data_in[208]&H_in[2256])^(data_in[209]&H_in[2257])^(data_in[210]&H_in[2258])^(data_in[211]&H_in[2259])^(data_in[212]&H_in[2260])^(data_in[213]&H_in[2261])^(data_in[214]&H_in[2262])^(data_in[215]&H_in[2263])^(data_in[216]&H_in[2264])^(data_in[217]&H_in[2265])^(data_in[218]&H_in[2266])^(data_in[219]&H_in[2267])^(data_in[220]&H_in[2268])^(data_in[221]&H_in[2269])^(data_in[222]&H_in[2270])^(data_in[223]&H_in[2271])^(data_in[224]&H_in[2272])^(data_in[225]&H_in[2273])^(data_in[226]&H_in[2274])^(data_in[227]&H_in[2275])^(data_in[228]&H_in[2276])^(data_in[229]&H_in[2277])^(data_in[230]&H_in[2278])^(data_in[231]&H_in[2279])^(data_in[232]&H_in[2280])^(data_in[233]&H_in[2281])^(data_in[234]&H_in[2282])^(data_in[235]&H_in[2283])^(data_in[236]&H_in[2284])^(data_in[237]&H_in[2285])^(data_in[238]&H_in[2286])^(data_in[239]&H_in[2287])^(data_in[240]&H_in[2288])^(data_in[241]&H_in[2289])^(data_in[242]&H_in[2290])^(data_in[243]&H_in[2291])^(data_in[244]&H_in[2292])^(data_in[245]&H_in[2293])^(data_in[246]&H_in[2294])^(data_in[247]&H_in[2295])^(data_in[248]&H_in[2296])^(data_in[249]&H_in[2297])^(data_in[250]&H_in[2298])^(data_in[251]&H_in[2299])^(data_in[252]&H_in[2300])^(data_in[253]&H_in[2301])^(data_in[254]&H_in[2302])^(data_in[255]&H_in[2303]);
         data_out[9]<=data_out[9]^(data_in[0]&H_in[2304])^(data_in[1]&H_in[2305])^(data_in[2]&H_in[2306])^(data_in[3]&H_in[2307])^(data_in[4]&H_in[2308])^(data_in[5]&H_in[2309])^(data_in[6]&H_in[2310])^(data_in[7]&H_in[2311])^(data_in[8]&H_in[2312])^(data_in[9]&H_in[2313])^(data_in[10]&H_in[2314])^(data_in[11]&H_in[2315])^(data_in[12]&H_in[2316])^(data_in[13]&H_in[2317])^(data_in[14]&H_in[2318])^(data_in[15]&H_in[2319])^(data_in[16]&H_in[2320])^(data_in[17]&H_in[2321])^(data_in[18]&H_in[2322])^(data_in[19]&H_in[2323])^(data_in[20]&H_in[2324])^(data_in[21]&H_in[2325])^(data_in[22]&H_in[2326])^(data_in[23]&H_in[2327])^(data_in[24]&H_in[2328])^(data_in[25]&H_in[2329])^(data_in[26]&H_in[2330])^(data_in[27]&H_in[2331])^(data_in[28]&H_in[2332])^(data_in[29]&H_in[2333])^(data_in[30]&H_in[2334])^(data_in[31]&H_in[2335])^(data_in[32]&H_in[2336])^(data_in[33]&H_in[2337])^(data_in[34]&H_in[2338])^(data_in[35]&H_in[2339])^(data_in[36]&H_in[2340])^(data_in[37]&H_in[2341])^(data_in[38]&H_in[2342])^(data_in[39]&H_in[2343])^(data_in[40]&H_in[2344])^(data_in[41]&H_in[2345])^(data_in[42]&H_in[2346])^(data_in[43]&H_in[2347])^(data_in[44]&H_in[2348])^(data_in[45]&H_in[2349])^(data_in[46]&H_in[2350])^(data_in[47]&H_in[2351])^(data_in[48]&H_in[2352])^(data_in[49]&H_in[2353])^(data_in[50]&H_in[2354])^(data_in[51]&H_in[2355])^(data_in[52]&H_in[2356])^(data_in[53]&H_in[2357])^(data_in[54]&H_in[2358])^(data_in[55]&H_in[2359])^(data_in[56]&H_in[2360])^(data_in[57]&H_in[2361])^(data_in[58]&H_in[2362])^(data_in[59]&H_in[2363])^(data_in[60]&H_in[2364])^(data_in[61]&H_in[2365])^(data_in[62]&H_in[2366])^(data_in[63]&H_in[2367])^(data_in[64]&H_in[2368])^(data_in[65]&H_in[2369])^(data_in[66]&H_in[2370])^(data_in[67]&H_in[2371])^(data_in[68]&H_in[2372])^(data_in[69]&H_in[2373])^(data_in[70]&H_in[2374])^(data_in[71]&H_in[2375])^(data_in[72]&H_in[2376])^(data_in[73]&H_in[2377])^(data_in[74]&H_in[2378])^(data_in[75]&H_in[2379])^(data_in[76]&H_in[2380])^(data_in[77]&H_in[2381])^(data_in[78]&H_in[2382])^(data_in[79]&H_in[2383])^(data_in[80]&H_in[2384])^(data_in[81]&H_in[2385])^(data_in[82]&H_in[2386])^(data_in[83]&H_in[2387])^(data_in[84]&H_in[2388])^(data_in[85]&H_in[2389])^(data_in[86]&H_in[2390])^(data_in[87]&H_in[2391])^(data_in[88]&H_in[2392])^(data_in[89]&H_in[2393])^(data_in[90]&H_in[2394])^(data_in[91]&H_in[2395])^(data_in[92]&H_in[2396])^(data_in[93]&H_in[2397])^(data_in[94]&H_in[2398])^(data_in[95]&H_in[2399])^(data_in[96]&H_in[2400])^(data_in[97]&H_in[2401])^(data_in[98]&H_in[2402])^(data_in[99]&H_in[2403])^(data_in[100]&H_in[2404])^(data_in[101]&H_in[2405])^(data_in[102]&H_in[2406])^(data_in[103]&H_in[2407])^(data_in[104]&H_in[2408])^(data_in[105]&H_in[2409])^(data_in[106]&H_in[2410])^(data_in[107]&H_in[2411])^(data_in[108]&H_in[2412])^(data_in[109]&H_in[2413])^(data_in[110]&H_in[2414])^(data_in[111]&H_in[2415])^(data_in[112]&H_in[2416])^(data_in[113]&H_in[2417])^(data_in[114]&H_in[2418])^(data_in[115]&H_in[2419])^(data_in[116]&H_in[2420])^(data_in[117]&H_in[2421])^(data_in[118]&H_in[2422])^(data_in[119]&H_in[2423])^(data_in[120]&H_in[2424])^(data_in[121]&H_in[2425])^(data_in[122]&H_in[2426])^(data_in[123]&H_in[2427])^(data_in[124]&H_in[2428])^(data_in[125]&H_in[2429])^(data_in[126]&H_in[2430])^(data_in[127]&H_in[2431])^(data_in[128]&H_in[2432])^(data_in[129]&H_in[2433])^(data_in[130]&H_in[2434])^(data_in[131]&H_in[2435])^(data_in[132]&H_in[2436])^(data_in[133]&H_in[2437])^(data_in[134]&H_in[2438])^(data_in[135]&H_in[2439])^(data_in[136]&H_in[2440])^(data_in[137]&H_in[2441])^(data_in[138]&H_in[2442])^(data_in[139]&H_in[2443])^(data_in[140]&H_in[2444])^(data_in[141]&H_in[2445])^(data_in[142]&H_in[2446])^(data_in[143]&H_in[2447])^(data_in[144]&H_in[2448])^(data_in[145]&H_in[2449])^(data_in[146]&H_in[2450])^(data_in[147]&H_in[2451])^(data_in[148]&H_in[2452])^(data_in[149]&H_in[2453])^(data_in[150]&H_in[2454])^(data_in[151]&H_in[2455])^(data_in[152]&H_in[2456])^(data_in[153]&H_in[2457])^(data_in[154]&H_in[2458])^(data_in[155]&H_in[2459])^(data_in[156]&H_in[2460])^(data_in[157]&H_in[2461])^(data_in[158]&H_in[2462])^(data_in[159]&H_in[2463])^(data_in[160]&H_in[2464])^(data_in[161]&H_in[2465])^(data_in[162]&H_in[2466])^(data_in[163]&H_in[2467])^(data_in[164]&H_in[2468])^(data_in[165]&H_in[2469])^(data_in[166]&H_in[2470])^(data_in[167]&H_in[2471])^(data_in[168]&H_in[2472])^(data_in[169]&H_in[2473])^(data_in[170]&H_in[2474])^(data_in[171]&H_in[2475])^(data_in[172]&H_in[2476])^(data_in[173]&H_in[2477])^(data_in[174]&H_in[2478])^(data_in[175]&H_in[2479])^(data_in[176]&H_in[2480])^(data_in[177]&H_in[2481])^(data_in[178]&H_in[2482])^(data_in[179]&H_in[2483])^(data_in[180]&H_in[2484])^(data_in[181]&H_in[2485])^(data_in[182]&H_in[2486])^(data_in[183]&H_in[2487])^(data_in[184]&H_in[2488])^(data_in[185]&H_in[2489])^(data_in[186]&H_in[2490])^(data_in[187]&H_in[2491])^(data_in[188]&H_in[2492])^(data_in[189]&H_in[2493])^(data_in[190]&H_in[2494])^(data_in[191]&H_in[2495])^(data_in[192]&H_in[2496])^(data_in[193]&H_in[2497])^(data_in[194]&H_in[2498])^(data_in[195]&H_in[2499])^(data_in[196]&H_in[2500])^(data_in[197]&H_in[2501])^(data_in[198]&H_in[2502])^(data_in[199]&H_in[2503])^(data_in[200]&H_in[2504])^(data_in[201]&H_in[2505])^(data_in[202]&H_in[2506])^(data_in[203]&H_in[2507])^(data_in[204]&H_in[2508])^(data_in[205]&H_in[2509])^(data_in[206]&H_in[2510])^(data_in[207]&H_in[2511])^(data_in[208]&H_in[2512])^(data_in[209]&H_in[2513])^(data_in[210]&H_in[2514])^(data_in[211]&H_in[2515])^(data_in[212]&H_in[2516])^(data_in[213]&H_in[2517])^(data_in[214]&H_in[2518])^(data_in[215]&H_in[2519])^(data_in[216]&H_in[2520])^(data_in[217]&H_in[2521])^(data_in[218]&H_in[2522])^(data_in[219]&H_in[2523])^(data_in[220]&H_in[2524])^(data_in[221]&H_in[2525])^(data_in[222]&H_in[2526])^(data_in[223]&H_in[2527])^(data_in[224]&H_in[2528])^(data_in[225]&H_in[2529])^(data_in[226]&H_in[2530])^(data_in[227]&H_in[2531])^(data_in[228]&H_in[2532])^(data_in[229]&H_in[2533])^(data_in[230]&H_in[2534])^(data_in[231]&H_in[2535])^(data_in[232]&H_in[2536])^(data_in[233]&H_in[2537])^(data_in[234]&H_in[2538])^(data_in[235]&H_in[2539])^(data_in[236]&H_in[2540])^(data_in[237]&H_in[2541])^(data_in[238]&H_in[2542])^(data_in[239]&H_in[2543])^(data_in[240]&H_in[2544])^(data_in[241]&H_in[2545])^(data_in[242]&H_in[2546])^(data_in[243]&H_in[2547])^(data_in[244]&H_in[2548])^(data_in[245]&H_in[2549])^(data_in[246]&H_in[2550])^(data_in[247]&H_in[2551])^(data_in[248]&H_in[2552])^(data_in[249]&H_in[2553])^(data_in[250]&H_in[2554])^(data_in[251]&H_in[2555])^(data_in[252]&H_in[2556])^(data_in[253]&H_in[2557])^(data_in[254]&H_in[2558])^(data_in[255]&H_in[2559]);
         data_out[10]<=data_out[10]^(data_in[0]&H_in[2560])^(data_in[1]&H_in[2561])^(data_in[2]&H_in[2562])^(data_in[3]&H_in[2563])^(data_in[4]&H_in[2564])^(data_in[5]&H_in[2565])^(data_in[6]&H_in[2566])^(data_in[7]&H_in[2567])^(data_in[8]&H_in[2568])^(data_in[9]&H_in[2569])^(data_in[10]&H_in[2570])^(data_in[11]&H_in[2571])^(data_in[12]&H_in[2572])^(data_in[13]&H_in[2573])^(data_in[14]&H_in[2574])^(data_in[15]&H_in[2575])^(data_in[16]&H_in[2576])^(data_in[17]&H_in[2577])^(data_in[18]&H_in[2578])^(data_in[19]&H_in[2579])^(data_in[20]&H_in[2580])^(data_in[21]&H_in[2581])^(data_in[22]&H_in[2582])^(data_in[23]&H_in[2583])^(data_in[24]&H_in[2584])^(data_in[25]&H_in[2585])^(data_in[26]&H_in[2586])^(data_in[27]&H_in[2587])^(data_in[28]&H_in[2588])^(data_in[29]&H_in[2589])^(data_in[30]&H_in[2590])^(data_in[31]&H_in[2591])^(data_in[32]&H_in[2592])^(data_in[33]&H_in[2593])^(data_in[34]&H_in[2594])^(data_in[35]&H_in[2595])^(data_in[36]&H_in[2596])^(data_in[37]&H_in[2597])^(data_in[38]&H_in[2598])^(data_in[39]&H_in[2599])^(data_in[40]&H_in[2600])^(data_in[41]&H_in[2601])^(data_in[42]&H_in[2602])^(data_in[43]&H_in[2603])^(data_in[44]&H_in[2604])^(data_in[45]&H_in[2605])^(data_in[46]&H_in[2606])^(data_in[47]&H_in[2607])^(data_in[48]&H_in[2608])^(data_in[49]&H_in[2609])^(data_in[50]&H_in[2610])^(data_in[51]&H_in[2611])^(data_in[52]&H_in[2612])^(data_in[53]&H_in[2613])^(data_in[54]&H_in[2614])^(data_in[55]&H_in[2615])^(data_in[56]&H_in[2616])^(data_in[57]&H_in[2617])^(data_in[58]&H_in[2618])^(data_in[59]&H_in[2619])^(data_in[60]&H_in[2620])^(data_in[61]&H_in[2621])^(data_in[62]&H_in[2622])^(data_in[63]&H_in[2623])^(data_in[64]&H_in[2624])^(data_in[65]&H_in[2625])^(data_in[66]&H_in[2626])^(data_in[67]&H_in[2627])^(data_in[68]&H_in[2628])^(data_in[69]&H_in[2629])^(data_in[70]&H_in[2630])^(data_in[71]&H_in[2631])^(data_in[72]&H_in[2632])^(data_in[73]&H_in[2633])^(data_in[74]&H_in[2634])^(data_in[75]&H_in[2635])^(data_in[76]&H_in[2636])^(data_in[77]&H_in[2637])^(data_in[78]&H_in[2638])^(data_in[79]&H_in[2639])^(data_in[80]&H_in[2640])^(data_in[81]&H_in[2641])^(data_in[82]&H_in[2642])^(data_in[83]&H_in[2643])^(data_in[84]&H_in[2644])^(data_in[85]&H_in[2645])^(data_in[86]&H_in[2646])^(data_in[87]&H_in[2647])^(data_in[88]&H_in[2648])^(data_in[89]&H_in[2649])^(data_in[90]&H_in[2650])^(data_in[91]&H_in[2651])^(data_in[92]&H_in[2652])^(data_in[93]&H_in[2653])^(data_in[94]&H_in[2654])^(data_in[95]&H_in[2655])^(data_in[96]&H_in[2656])^(data_in[97]&H_in[2657])^(data_in[98]&H_in[2658])^(data_in[99]&H_in[2659])^(data_in[100]&H_in[2660])^(data_in[101]&H_in[2661])^(data_in[102]&H_in[2662])^(data_in[103]&H_in[2663])^(data_in[104]&H_in[2664])^(data_in[105]&H_in[2665])^(data_in[106]&H_in[2666])^(data_in[107]&H_in[2667])^(data_in[108]&H_in[2668])^(data_in[109]&H_in[2669])^(data_in[110]&H_in[2670])^(data_in[111]&H_in[2671])^(data_in[112]&H_in[2672])^(data_in[113]&H_in[2673])^(data_in[114]&H_in[2674])^(data_in[115]&H_in[2675])^(data_in[116]&H_in[2676])^(data_in[117]&H_in[2677])^(data_in[118]&H_in[2678])^(data_in[119]&H_in[2679])^(data_in[120]&H_in[2680])^(data_in[121]&H_in[2681])^(data_in[122]&H_in[2682])^(data_in[123]&H_in[2683])^(data_in[124]&H_in[2684])^(data_in[125]&H_in[2685])^(data_in[126]&H_in[2686])^(data_in[127]&H_in[2687])^(data_in[128]&H_in[2688])^(data_in[129]&H_in[2689])^(data_in[130]&H_in[2690])^(data_in[131]&H_in[2691])^(data_in[132]&H_in[2692])^(data_in[133]&H_in[2693])^(data_in[134]&H_in[2694])^(data_in[135]&H_in[2695])^(data_in[136]&H_in[2696])^(data_in[137]&H_in[2697])^(data_in[138]&H_in[2698])^(data_in[139]&H_in[2699])^(data_in[140]&H_in[2700])^(data_in[141]&H_in[2701])^(data_in[142]&H_in[2702])^(data_in[143]&H_in[2703])^(data_in[144]&H_in[2704])^(data_in[145]&H_in[2705])^(data_in[146]&H_in[2706])^(data_in[147]&H_in[2707])^(data_in[148]&H_in[2708])^(data_in[149]&H_in[2709])^(data_in[150]&H_in[2710])^(data_in[151]&H_in[2711])^(data_in[152]&H_in[2712])^(data_in[153]&H_in[2713])^(data_in[154]&H_in[2714])^(data_in[155]&H_in[2715])^(data_in[156]&H_in[2716])^(data_in[157]&H_in[2717])^(data_in[158]&H_in[2718])^(data_in[159]&H_in[2719])^(data_in[160]&H_in[2720])^(data_in[161]&H_in[2721])^(data_in[162]&H_in[2722])^(data_in[163]&H_in[2723])^(data_in[164]&H_in[2724])^(data_in[165]&H_in[2725])^(data_in[166]&H_in[2726])^(data_in[167]&H_in[2727])^(data_in[168]&H_in[2728])^(data_in[169]&H_in[2729])^(data_in[170]&H_in[2730])^(data_in[171]&H_in[2731])^(data_in[172]&H_in[2732])^(data_in[173]&H_in[2733])^(data_in[174]&H_in[2734])^(data_in[175]&H_in[2735])^(data_in[176]&H_in[2736])^(data_in[177]&H_in[2737])^(data_in[178]&H_in[2738])^(data_in[179]&H_in[2739])^(data_in[180]&H_in[2740])^(data_in[181]&H_in[2741])^(data_in[182]&H_in[2742])^(data_in[183]&H_in[2743])^(data_in[184]&H_in[2744])^(data_in[185]&H_in[2745])^(data_in[186]&H_in[2746])^(data_in[187]&H_in[2747])^(data_in[188]&H_in[2748])^(data_in[189]&H_in[2749])^(data_in[190]&H_in[2750])^(data_in[191]&H_in[2751])^(data_in[192]&H_in[2752])^(data_in[193]&H_in[2753])^(data_in[194]&H_in[2754])^(data_in[195]&H_in[2755])^(data_in[196]&H_in[2756])^(data_in[197]&H_in[2757])^(data_in[198]&H_in[2758])^(data_in[199]&H_in[2759])^(data_in[200]&H_in[2760])^(data_in[201]&H_in[2761])^(data_in[202]&H_in[2762])^(data_in[203]&H_in[2763])^(data_in[204]&H_in[2764])^(data_in[205]&H_in[2765])^(data_in[206]&H_in[2766])^(data_in[207]&H_in[2767])^(data_in[208]&H_in[2768])^(data_in[209]&H_in[2769])^(data_in[210]&H_in[2770])^(data_in[211]&H_in[2771])^(data_in[212]&H_in[2772])^(data_in[213]&H_in[2773])^(data_in[214]&H_in[2774])^(data_in[215]&H_in[2775])^(data_in[216]&H_in[2776])^(data_in[217]&H_in[2777])^(data_in[218]&H_in[2778])^(data_in[219]&H_in[2779])^(data_in[220]&H_in[2780])^(data_in[221]&H_in[2781])^(data_in[222]&H_in[2782])^(data_in[223]&H_in[2783])^(data_in[224]&H_in[2784])^(data_in[225]&H_in[2785])^(data_in[226]&H_in[2786])^(data_in[227]&H_in[2787])^(data_in[228]&H_in[2788])^(data_in[229]&H_in[2789])^(data_in[230]&H_in[2790])^(data_in[231]&H_in[2791])^(data_in[232]&H_in[2792])^(data_in[233]&H_in[2793])^(data_in[234]&H_in[2794])^(data_in[235]&H_in[2795])^(data_in[236]&H_in[2796])^(data_in[237]&H_in[2797])^(data_in[238]&H_in[2798])^(data_in[239]&H_in[2799])^(data_in[240]&H_in[2800])^(data_in[241]&H_in[2801])^(data_in[242]&H_in[2802])^(data_in[243]&H_in[2803])^(data_in[244]&H_in[2804])^(data_in[245]&H_in[2805])^(data_in[246]&H_in[2806])^(data_in[247]&H_in[2807])^(data_in[248]&H_in[2808])^(data_in[249]&H_in[2809])^(data_in[250]&H_in[2810])^(data_in[251]&H_in[2811])^(data_in[252]&H_in[2812])^(data_in[253]&H_in[2813])^(data_in[254]&H_in[2814])^(data_in[255]&H_in[2815]);
         data_out[11]<=data_out[11]^(data_in[0]&H_in[2816])^(data_in[1]&H_in[2817])^(data_in[2]&H_in[2818])^(data_in[3]&H_in[2819])^(data_in[4]&H_in[2820])^(data_in[5]&H_in[2821])^(data_in[6]&H_in[2822])^(data_in[7]&H_in[2823])^(data_in[8]&H_in[2824])^(data_in[9]&H_in[2825])^(data_in[10]&H_in[2826])^(data_in[11]&H_in[2827])^(data_in[12]&H_in[2828])^(data_in[13]&H_in[2829])^(data_in[14]&H_in[2830])^(data_in[15]&H_in[2831])^(data_in[16]&H_in[2832])^(data_in[17]&H_in[2833])^(data_in[18]&H_in[2834])^(data_in[19]&H_in[2835])^(data_in[20]&H_in[2836])^(data_in[21]&H_in[2837])^(data_in[22]&H_in[2838])^(data_in[23]&H_in[2839])^(data_in[24]&H_in[2840])^(data_in[25]&H_in[2841])^(data_in[26]&H_in[2842])^(data_in[27]&H_in[2843])^(data_in[28]&H_in[2844])^(data_in[29]&H_in[2845])^(data_in[30]&H_in[2846])^(data_in[31]&H_in[2847])^(data_in[32]&H_in[2848])^(data_in[33]&H_in[2849])^(data_in[34]&H_in[2850])^(data_in[35]&H_in[2851])^(data_in[36]&H_in[2852])^(data_in[37]&H_in[2853])^(data_in[38]&H_in[2854])^(data_in[39]&H_in[2855])^(data_in[40]&H_in[2856])^(data_in[41]&H_in[2857])^(data_in[42]&H_in[2858])^(data_in[43]&H_in[2859])^(data_in[44]&H_in[2860])^(data_in[45]&H_in[2861])^(data_in[46]&H_in[2862])^(data_in[47]&H_in[2863])^(data_in[48]&H_in[2864])^(data_in[49]&H_in[2865])^(data_in[50]&H_in[2866])^(data_in[51]&H_in[2867])^(data_in[52]&H_in[2868])^(data_in[53]&H_in[2869])^(data_in[54]&H_in[2870])^(data_in[55]&H_in[2871])^(data_in[56]&H_in[2872])^(data_in[57]&H_in[2873])^(data_in[58]&H_in[2874])^(data_in[59]&H_in[2875])^(data_in[60]&H_in[2876])^(data_in[61]&H_in[2877])^(data_in[62]&H_in[2878])^(data_in[63]&H_in[2879])^(data_in[64]&H_in[2880])^(data_in[65]&H_in[2881])^(data_in[66]&H_in[2882])^(data_in[67]&H_in[2883])^(data_in[68]&H_in[2884])^(data_in[69]&H_in[2885])^(data_in[70]&H_in[2886])^(data_in[71]&H_in[2887])^(data_in[72]&H_in[2888])^(data_in[73]&H_in[2889])^(data_in[74]&H_in[2890])^(data_in[75]&H_in[2891])^(data_in[76]&H_in[2892])^(data_in[77]&H_in[2893])^(data_in[78]&H_in[2894])^(data_in[79]&H_in[2895])^(data_in[80]&H_in[2896])^(data_in[81]&H_in[2897])^(data_in[82]&H_in[2898])^(data_in[83]&H_in[2899])^(data_in[84]&H_in[2900])^(data_in[85]&H_in[2901])^(data_in[86]&H_in[2902])^(data_in[87]&H_in[2903])^(data_in[88]&H_in[2904])^(data_in[89]&H_in[2905])^(data_in[90]&H_in[2906])^(data_in[91]&H_in[2907])^(data_in[92]&H_in[2908])^(data_in[93]&H_in[2909])^(data_in[94]&H_in[2910])^(data_in[95]&H_in[2911])^(data_in[96]&H_in[2912])^(data_in[97]&H_in[2913])^(data_in[98]&H_in[2914])^(data_in[99]&H_in[2915])^(data_in[100]&H_in[2916])^(data_in[101]&H_in[2917])^(data_in[102]&H_in[2918])^(data_in[103]&H_in[2919])^(data_in[104]&H_in[2920])^(data_in[105]&H_in[2921])^(data_in[106]&H_in[2922])^(data_in[107]&H_in[2923])^(data_in[108]&H_in[2924])^(data_in[109]&H_in[2925])^(data_in[110]&H_in[2926])^(data_in[111]&H_in[2927])^(data_in[112]&H_in[2928])^(data_in[113]&H_in[2929])^(data_in[114]&H_in[2930])^(data_in[115]&H_in[2931])^(data_in[116]&H_in[2932])^(data_in[117]&H_in[2933])^(data_in[118]&H_in[2934])^(data_in[119]&H_in[2935])^(data_in[120]&H_in[2936])^(data_in[121]&H_in[2937])^(data_in[122]&H_in[2938])^(data_in[123]&H_in[2939])^(data_in[124]&H_in[2940])^(data_in[125]&H_in[2941])^(data_in[126]&H_in[2942])^(data_in[127]&H_in[2943])^(data_in[128]&H_in[2944])^(data_in[129]&H_in[2945])^(data_in[130]&H_in[2946])^(data_in[131]&H_in[2947])^(data_in[132]&H_in[2948])^(data_in[133]&H_in[2949])^(data_in[134]&H_in[2950])^(data_in[135]&H_in[2951])^(data_in[136]&H_in[2952])^(data_in[137]&H_in[2953])^(data_in[138]&H_in[2954])^(data_in[139]&H_in[2955])^(data_in[140]&H_in[2956])^(data_in[141]&H_in[2957])^(data_in[142]&H_in[2958])^(data_in[143]&H_in[2959])^(data_in[144]&H_in[2960])^(data_in[145]&H_in[2961])^(data_in[146]&H_in[2962])^(data_in[147]&H_in[2963])^(data_in[148]&H_in[2964])^(data_in[149]&H_in[2965])^(data_in[150]&H_in[2966])^(data_in[151]&H_in[2967])^(data_in[152]&H_in[2968])^(data_in[153]&H_in[2969])^(data_in[154]&H_in[2970])^(data_in[155]&H_in[2971])^(data_in[156]&H_in[2972])^(data_in[157]&H_in[2973])^(data_in[158]&H_in[2974])^(data_in[159]&H_in[2975])^(data_in[160]&H_in[2976])^(data_in[161]&H_in[2977])^(data_in[162]&H_in[2978])^(data_in[163]&H_in[2979])^(data_in[164]&H_in[2980])^(data_in[165]&H_in[2981])^(data_in[166]&H_in[2982])^(data_in[167]&H_in[2983])^(data_in[168]&H_in[2984])^(data_in[169]&H_in[2985])^(data_in[170]&H_in[2986])^(data_in[171]&H_in[2987])^(data_in[172]&H_in[2988])^(data_in[173]&H_in[2989])^(data_in[174]&H_in[2990])^(data_in[175]&H_in[2991])^(data_in[176]&H_in[2992])^(data_in[177]&H_in[2993])^(data_in[178]&H_in[2994])^(data_in[179]&H_in[2995])^(data_in[180]&H_in[2996])^(data_in[181]&H_in[2997])^(data_in[182]&H_in[2998])^(data_in[183]&H_in[2999])^(data_in[184]&H_in[3000])^(data_in[185]&H_in[3001])^(data_in[186]&H_in[3002])^(data_in[187]&H_in[3003])^(data_in[188]&H_in[3004])^(data_in[189]&H_in[3005])^(data_in[190]&H_in[3006])^(data_in[191]&H_in[3007])^(data_in[192]&H_in[3008])^(data_in[193]&H_in[3009])^(data_in[194]&H_in[3010])^(data_in[195]&H_in[3011])^(data_in[196]&H_in[3012])^(data_in[197]&H_in[3013])^(data_in[198]&H_in[3014])^(data_in[199]&H_in[3015])^(data_in[200]&H_in[3016])^(data_in[201]&H_in[3017])^(data_in[202]&H_in[3018])^(data_in[203]&H_in[3019])^(data_in[204]&H_in[3020])^(data_in[205]&H_in[3021])^(data_in[206]&H_in[3022])^(data_in[207]&H_in[3023])^(data_in[208]&H_in[3024])^(data_in[209]&H_in[3025])^(data_in[210]&H_in[3026])^(data_in[211]&H_in[3027])^(data_in[212]&H_in[3028])^(data_in[213]&H_in[3029])^(data_in[214]&H_in[3030])^(data_in[215]&H_in[3031])^(data_in[216]&H_in[3032])^(data_in[217]&H_in[3033])^(data_in[218]&H_in[3034])^(data_in[219]&H_in[3035])^(data_in[220]&H_in[3036])^(data_in[221]&H_in[3037])^(data_in[222]&H_in[3038])^(data_in[223]&H_in[3039])^(data_in[224]&H_in[3040])^(data_in[225]&H_in[3041])^(data_in[226]&H_in[3042])^(data_in[227]&H_in[3043])^(data_in[228]&H_in[3044])^(data_in[229]&H_in[3045])^(data_in[230]&H_in[3046])^(data_in[231]&H_in[3047])^(data_in[232]&H_in[3048])^(data_in[233]&H_in[3049])^(data_in[234]&H_in[3050])^(data_in[235]&H_in[3051])^(data_in[236]&H_in[3052])^(data_in[237]&H_in[3053])^(data_in[238]&H_in[3054])^(data_in[239]&H_in[3055])^(data_in[240]&H_in[3056])^(data_in[241]&H_in[3057])^(data_in[242]&H_in[3058])^(data_in[243]&H_in[3059])^(data_in[244]&H_in[3060])^(data_in[245]&H_in[3061])^(data_in[246]&H_in[3062])^(data_in[247]&H_in[3063])^(data_in[248]&H_in[3064])^(data_in[249]&H_in[3065])^(data_in[250]&H_in[3066])^(data_in[251]&H_in[3067])^(data_in[252]&H_in[3068])^(data_in[253]&H_in[3069])^(data_in[254]&H_in[3070])^(data_in[255]&H_in[3071]);
         data_out[12]<=data_out[12]^(data_in[0]&H_in[3072])^(data_in[1]&H_in[3073])^(data_in[2]&H_in[3074])^(data_in[3]&H_in[3075])^(data_in[4]&H_in[3076])^(data_in[5]&H_in[3077])^(data_in[6]&H_in[3078])^(data_in[7]&H_in[3079])^(data_in[8]&H_in[3080])^(data_in[9]&H_in[3081])^(data_in[10]&H_in[3082])^(data_in[11]&H_in[3083])^(data_in[12]&H_in[3084])^(data_in[13]&H_in[3085])^(data_in[14]&H_in[3086])^(data_in[15]&H_in[3087])^(data_in[16]&H_in[3088])^(data_in[17]&H_in[3089])^(data_in[18]&H_in[3090])^(data_in[19]&H_in[3091])^(data_in[20]&H_in[3092])^(data_in[21]&H_in[3093])^(data_in[22]&H_in[3094])^(data_in[23]&H_in[3095])^(data_in[24]&H_in[3096])^(data_in[25]&H_in[3097])^(data_in[26]&H_in[3098])^(data_in[27]&H_in[3099])^(data_in[28]&H_in[3100])^(data_in[29]&H_in[3101])^(data_in[30]&H_in[3102])^(data_in[31]&H_in[3103])^(data_in[32]&H_in[3104])^(data_in[33]&H_in[3105])^(data_in[34]&H_in[3106])^(data_in[35]&H_in[3107])^(data_in[36]&H_in[3108])^(data_in[37]&H_in[3109])^(data_in[38]&H_in[3110])^(data_in[39]&H_in[3111])^(data_in[40]&H_in[3112])^(data_in[41]&H_in[3113])^(data_in[42]&H_in[3114])^(data_in[43]&H_in[3115])^(data_in[44]&H_in[3116])^(data_in[45]&H_in[3117])^(data_in[46]&H_in[3118])^(data_in[47]&H_in[3119])^(data_in[48]&H_in[3120])^(data_in[49]&H_in[3121])^(data_in[50]&H_in[3122])^(data_in[51]&H_in[3123])^(data_in[52]&H_in[3124])^(data_in[53]&H_in[3125])^(data_in[54]&H_in[3126])^(data_in[55]&H_in[3127])^(data_in[56]&H_in[3128])^(data_in[57]&H_in[3129])^(data_in[58]&H_in[3130])^(data_in[59]&H_in[3131])^(data_in[60]&H_in[3132])^(data_in[61]&H_in[3133])^(data_in[62]&H_in[3134])^(data_in[63]&H_in[3135])^(data_in[64]&H_in[3136])^(data_in[65]&H_in[3137])^(data_in[66]&H_in[3138])^(data_in[67]&H_in[3139])^(data_in[68]&H_in[3140])^(data_in[69]&H_in[3141])^(data_in[70]&H_in[3142])^(data_in[71]&H_in[3143])^(data_in[72]&H_in[3144])^(data_in[73]&H_in[3145])^(data_in[74]&H_in[3146])^(data_in[75]&H_in[3147])^(data_in[76]&H_in[3148])^(data_in[77]&H_in[3149])^(data_in[78]&H_in[3150])^(data_in[79]&H_in[3151])^(data_in[80]&H_in[3152])^(data_in[81]&H_in[3153])^(data_in[82]&H_in[3154])^(data_in[83]&H_in[3155])^(data_in[84]&H_in[3156])^(data_in[85]&H_in[3157])^(data_in[86]&H_in[3158])^(data_in[87]&H_in[3159])^(data_in[88]&H_in[3160])^(data_in[89]&H_in[3161])^(data_in[90]&H_in[3162])^(data_in[91]&H_in[3163])^(data_in[92]&H_in[3164])^(data_in[93]&H_in[3165])^(data_in[94]&H_in[3166])^(data_in[95]&H_in[3167])^(data_in[96]&H_in[3168])^(data_in[97]&H_in[3169])^(data_in[98]&H_in[3170])^(data_in[99]&H_in[3171])^(data_in[100]&H_in[3172])^(data_in[101]&H_in[3173])^(data_in[102]&H_in[3174])^(data_in[103]&H_in[3175])^(data_in[104]&H_in[3176])^(data_in[105]&H_in[3177])^(data_in[106]&H_in[3178])^(data_in[107]&H_in[3179])^(data_in[108]&H_in[3180])^(data_in[109]&H_in[3181])^(data_in[110]&H_in[3182])^(data_in[111]&H_in[3183])^(data_in[112]&H_in[3184])^(data_in[113]&H_in[3185])^(data_in[114]&H_in[3186])^(data_in[115]&H_in[3187])^(data_in[116]&H_in[3188])^(data_in[117]&H_in[3189])^(data_in[118]&H_in[3190])^(data_in[119]&H_in[3191])^(data_in[120]&H_in[3192])^(data_in[121]&H_in[3193])^(data_in[122]&H_in[3194])^(data_in[123]&H_in[3195])^(data_in[124]&H_in[3196])^(data_in[125]&H_in[3197])^(data_in[126]&H_in[3198])^(data_in[127]&H_in[3199])^(data_in[128]&H_in[3200])^(data_in[129]&H_in[3201])^(data_in[130]&H_in[3202])^(data_in[131]&H_in[3203])^(data_in[132]&H_in[3204])^(data_in[133]&H_in[3205])^(data_in[134]&H_in[3206])^(data_in[135]&H_in[3207])^(data_in[136]&H_in[3208])^(data_in[137]&H_in[3209])^(data_in[138]&H_in[3210])^(data_in[139]&H_in[3211])^(data_in[140]&H_in[3212])^(data_in[141]&H_in[3213])^(data_in[142]&H_in[3214])^(data_in[143]&H_in[3215])^(data_in[144]&H_in[3216])^(data_in[145]&H_in[3217])^(data_in[146]&H_in[3218])^(data_in[147]&H_in[3219])^(data_in[148]&H_in[3220])^(data_in[149]&H_in[3221])^(data_in[150]&H_in[3222])^(data_in[151]&H_in[3223])^(data_in[152]&H_in[3224])^(data_in[153]&H_in[3225])^(data_in[154]&H_in[3226])^(data_in[155]&H_in[3227])^(data_in[156]&H_in[3228])^(data_in[157]&H_in[3229])^(data_in[158]&H_in[3230])^(data_in[159]&H_in[3231])^(data_in[160]&H_in[3232])^(data_in[161]&H_in[3233])^(data_in[162]&H_in[3234])^(data_in[163]&H_in[3235])^(data_in[164]&H_in[3236])^(data_in[165]&H_in[3237])^(data_in[166]&H_in[3238])^(data_in[167]&H_in[3239])^(data_in[168]&H_in[3240])^(data_in[169]&H_in[3241])^(data_in[170]&H_in[3242])^(data_in[171]&H_in[3243])^(data_in[172]&H_in[3244])^(data_in[173]&H_in[3245])^(data_in[174]&H_in[3246])^(data_in[175]&H_in[3247])^(data_in[176]&H_in[3248])^(data_in[177]&H_in[3249])^(data_in[178]&H_in[3250])^(data_in[179]&H_in[3251])^(data_in[180]&H_in[3252])^(data_in[181]&H_in[3253])^(data_in[182]&H_in[3254])^(data_in[183]&H_in[3255])^(data_in[184]&H_in[3256])^(data_in[185]&H_in[3257])^(data_in[186]&H_in[3258])^(data_in[187]&H_in[3259])^(data_in[188]&H_in[3260])^(data_in[189]&H_in[3261])^(data_in[190]&H_in[3262])^(data_in[191]&H_in[3263])^(data_in[192]&H_in[3264])^(data_in[193]&H_in[3265])^(data_in[194]&H_in[3266])^(data_in[195]&H_in[3267])^(data_in[196]&H_in[3268])^(data_in[197]&H_in[3269])^(data_in[198]&H_in[3270])^(data_in[199]&H_in[3271])^(data_in[200]&H_in[3272])^(data_in[201]&H_in[3273])^(data_in[202]&H_in[3274])^(data_in[203]&H_in[3275])^(data_in[204]&H_in[3276])^(data_in[205]&H_in[3277])^(data_in[206]&H_in[3278])^(data_in[207]&H_in[3279])^(data_in[208]&H_in[3280])^(data_in[209]&H_in[3281])^(data_in[210]&H_in[3282])^(data_in[211]&H_in[3283])^(data_in[212]&H_in[3284])^(data_in[213]&H_in[3285])^(data_in[214]&H_in[3286])^(data_in[215]&H_in[3287])^(data_in[216]&H_in[3288])^(data_in[217]&H_in[3289])^(data_in[218]&H_in[3290])^(data_in[219]&H_in[3291])^(data_in[220]&H_in[3292])^(data_in[221]&H_in[3293])^(data_in[222]&H_in[3294])^(data_in[223]&H_in[3295])^(data_in[224]&H_in[3296])^(data_in[225]&H_in[3297])^(data_in[226]&H_in[3298])^(data_in[227]&H_in[3299])^(data_in[228]&H_in[3300])^(data_in[229]&H_in[3301])^(data_in[230]&H_in[3302])^(data_in[231]&H_in[3303])^(data_in[232]&H_in[3304])^(data_in[233]&H_in[3305])^(data_in[234]&H_in[3306])^(data_in[235]&H_in[3307])^(data_in[236]&H_in[3308])^(data_in[237]&H_in[3309])^(data_in[238]&H_in[3310])^(data_in[239]&H_in[3311])^(data_in[240]&H_in[3312])^(data_in[241]&H_in[3313])^(data_in[242]&H_in[3314])^(data_in[243]&H_in[3315])^(data_in[244]&H_in[3316])^(data_in[245]&H_in[3317])^(data_in[246]&H_in[3318])^(data_in[247]&H_in[3319])^(data_in[248]&H_in[3320])^(data_in[249]&H_in[3321])^(data_in[250]&H_in[3322])^(data_in[251]&H_in[3323])^(data_in[252]&H_in[3324])^(data_in[253]&H_in[3325])^(data_in[254]&H_in[3326])^(data_in[255]&H_in[3327]);
         data_out[13]<=data_out[13]^(data_in[0]&H_in[3328])^(data_in[1]&H_in[3329])^(data_in[2]&H_in[3330])^(data_in[3]&H_in[3331])^(data_in[4]&H_in[3332])^(data_in[5]&H_in[3333])^(data_in[6]&H_in[3334])^(data_in[7]&H_in[3335])^(data_in[8]&H_in[3336])^(data_in[9]&H_in[3337])^(data_in[10]&H_in[3338])^(data_in[11]&H_in[3339])^(data_in[12]&H_in[3340])^(data_in[13]&H_in[3341])^(data_in[14]&H_in[3342])^(data_in[15]&H_in[3343])^(data_in[16]&H_in[3344])^(data_in[17]&H_in[3345])^(data_in[18]&H_in[3346])^(data_in[19]&H_in[3347])^(data_in[20]&H_in[3348])^(data_in[21]&H_in[3349])^(data_in[22]&H_in[3350])^(data_in[23]&H_in[3351])^(data_in[24]&H_in[3352])^(data_in[25]&H_in[3353])^(data_in[26]&H_in[3354])^(data_in[27]&H_in[3355])^(data_in[28]&H_in[3356])^(data_in[29]&H_in[3357])^(data_in[30]&H_in[3358])^(data_in[31]&H_in[3359])^(data_in[32]&H_in[3360])^(data_in[33]&H_in[3361])^(data_in[34]&H_in[3362])^(data_in[35]&H_in[3363])^(data_in[36]&H_in[3364])^(data_in[37]&H_in[3365])^(data_in[38]&H_in[3366])^(data_in[39]&H_in[3367])^(data_in[40]&H_in[3368])^(data_in[41]&H_in[3369])^(data_in[42]&H_in[3370])^(data_in[43]&H_in[3371])^(data_in[44]&H_in[3372])^(data_in[45]&H_in[3373])^(data_in[46]&H_in[3374])^(data_in[47]&H_in[3375])^(data_in[48]&H_in[3376])^(data_in[49]&H_in[3377])^(data_in[50]&H_in[3378])^(data_in[51]&H_in[3379])^(data_in[52]&H_in[3380])^(data_in[53]&H_in[3381])^(data_in[54]&H_in[3382])^(data_in[55]&H_in[3383])^(data_in[56]&H_in[3384])^(data_in[57]&H_in[3385])^(data_in[58]&H_in[3386])^(data_in[59]&H_in[3387])^(data_in[60]&H_in[3388])^(data_in[61]&H_in[3389])^(data_in[62]&H_in[3390])^(data_in[63]&H_in[3391])^(data_in[64]&H_in[3392])^(data_in[65]&H_in[3393])^(data_in[66]&H_in[3394])^(data_in[67]&H_in[3395])^(data_in[68]&H_in[3396])^(data_in[69]&H_in[3397])^(data_in[70]&H_in[3398])^(data_in[71]&H_in[3399])^(data_in[72]&H_in[3400])^(data_in[73]&H_in[3401])^(data_in[74]&H_in[3402])^(data_in[75]&H_in[3403])^(data_in[76]&H_in[3404])^(data_in[77]&H_in[3405])^(data_in[78]&H_in[3406])^(data_in[79]&H_in[3407])^(data_in[80]&H_in[3408])^(data_in[81]&H_in[3409])^(data_in[82]&H_in[3410])^(data_in[83]&H_in[3411])^(data_in[84]&H_in[3412])^(data_in[85]&H_in[3413])^(data_in[86]&H_in[3414])^(data_in[87]&H_in[3415])^(data_in[88]&H_in[3416])^(data_in[89]&H_in[3417])^(data_in[90]&H_in[3418])^(data_in[91]&H_in[3419])^(data_in[92]&H_in[3420])^(data_in[93]&H_in[3421])^(data_in[94]&H_in[3422])^(data_in[95]&H_in[3423])^(data_in[96]&H_in[3424])^(data_in[97]&H_in[3425])^(data_in[98]&H_in[3426])^(data_in[99]&H_in[3427])^(data_in[100]&H_in[3428])^(data_in[101]&H_in[3429])^(data_in[102]&H_in[3430])^(data_in[103]&H_in[3431])^(data_in[104]&H_in[3432])^(data_in[105]&H_in[3433])^(data_in[106]&H_in[3434])^(data_in[107]&H_in[3435])^(data_in[108]&H_in[3436])^(data_in[109]&H_in[3437])^(data_in[110]&H_in[3438])^(data_in[111]&H_in[3439])^(data_in[112]&H_in[3440])^(data_in[113]&H_in[3441])^(data_in[114]&H_in[3442])^(data_in[115]&H_in[3443])^(data_in[116]&H_in[3444])^(data_in[117]&H_in[3445])^(data_in[118]&H_in[3446])^(data_in[119]&H_in[3447])^(data_in[120]&H_in[3448])^(data_in[121]&H_in[3449])^(data_in[122]&H_in[3450])^(data_in[123]&H_in[3451])^(data_in[124]&H_in[3452])^(data_in[125]&H_in[3453])^(data_in[126]&H_in[3454])^(data_in[127]&H_in[3455])^(data_in[128]&H_in[3456])^(data_in[129]&H_in[3457])^(data_in[130]&H_in[3458])^(data_in[131]&H_in[3459])^(data_in[132]&H_in[3460])^(data_in[133]&H_in[3461])^(data_in[134]&H_in[3462])^(data_in[135]&H_in[3463])^(data_in[136]&H_in[3464])^(data_in[137]&H_in[3465])^(data_in[138]&H_in[3466])^(data_in[139]&H_in[3467])^(data_in[140]&H_in[3468])^(data_in[141]&H_in[3469])^(data_in[142]&H_in[3470])^(data_in[143]&H_in[3471])^(data_in[144]&H_in[3472])^(data_in[145]&H_in[3473])^(data_in[146]&H_in[3474])^(data_in[147]&H_in[3475])^(data_in[148]&H_in[3476])^(data_in[149]&H_in[3477])^(data_in[150]&H_in[3478])^(data_in[151]&H_in[3479])^(data_in[152]&H_in[3480])^(data_in[153]&H_in[3481])^(data_in[154]&H_in[3482])^(data_in[155]&H_in[3483])^(data_in[156]&H_in[3484])^(data_in[157]&H_in[3485])^(data_in[158]&H_in[3486])^(data_in[159]&H_in[3487])^(data_in[160]&H_in[3488])^(data_in[161]&H_in[3489])^(data_in[162]&H_in[3490])^(data_in[163]&H_in[3491])^(data_in[164]&H_in[3492])^(data_in[165]&H_in[3493])^(data_in[166]&H_in[3494])^(data_in[167]&H_in[3495])^(data_in[168]&H_in[3496])^(data_in[169]&H_in[3497])^(data_in[170]&H_in[3498])^(data_in[171]&H_in[3499])^(data_in[172]&H_in[3500])^(data_in[173]&H_in[3501])^(data_in[174]&H_in[3502])^(data_in[175]&H_in[3503])^(data_in[176]&H_in[3504])^(data_in[177]&H_in[3505])^(data_in[178]&H_in[3506])^(data_in[179]&H_in[3507])^(data_in[180]&H_in[3508])^(data_in[181]&H_in[3509])^(data_in[182]&H_in[3510])^(data_in[183]&H_in[3511])^(data_in[184]&H_in[3512])^(data_in[185]&H_in[3513])^(data_in[186]&H_in[3514])^(data_in[187]&H_in[3515])^(data_in[188]&H_in[3516])^(data_in[189]&H_in[3517])^(data_in[190]&H_in[3518])^(data_in[191]&H_in[3519])^(data_in[192]&H_in[3520])^(data_in[193]&H_in[3521])^(data_in[194]&H_in[3522])^(data_in[195]&H_in[3523])^(data_in[196]&H_in[3524])^(data_in[197]&H_in[3525])^(data_in[198]&H_in[3526])^(data_in[199]&H_in[3527])^(data_in[200]&H_in[3528])^(data_in[201]&H_in[3529])^(data_in[202]&H_in[3530])^(data_in[203]&H_in[3531])^(data_in[204]&H_in[3532])^(data_in[205]&H_in[3533])^(data_in[206]&H_in[3534])^(data_in[207]&H_in[3535])^(data_in[208]&H_in[3536])^(data_in[209]&H_in[3537])^(data_in[210]&H_in[3538])^(data_in[211]&H_in[3539])^(data_in[212]&H_in[3540])^(data_in[213]&H_in[3541])^(data_in[214]&H_in[3542])^(data_in[215]&H_in[3543])^(data_in[216]&H_in[3544])^(data_in[217]&H_in[3545])^(data_in[218]&H_in[3546])^(data_in[219]&H_in[3547])^(data_in[220]&H_in[3548])^(data_in[221]&H_in[3549])^(data_in[222]&H_in[3550])^(data_in[223]&H_in[3551])^(data_in[224]&H_in[3552])^(data_in[225]&H_in[3553])^(data_in[226]&H_in[3554])^(data_in[227]&H_in[3555])^(data_in[228]&H_in[3556])^(data_in[229]&H_in[3557])^(data_in[230]&H_in[3558])^(data_in[231]&H_in[3559])^(data_in[232]&H_in[3560])^(data_in[233]&H_in[3561])^(data_in[234]&H_in[3562])^(data_in[235]&H_in[3563])^(data_in[236]&H_in[3564])^(data_in[237]&H_in[3565])^(data_in[238]&H_in[3566])^(data_in[239]&H_in[3567])^(data_in[240]&H_in[3568])^(data_in[241]&H_in[3569])^(data_in[242]&H_in[3570])^(data_in[243]&H_in[3571])^(data_in[244]&H_in[3572])^(data_in[245]&H_in[3573])^(data_in[246]&H_in[3574])^(data_in[247]&H_in[3575])^(data_in[248]&H_in[3576])^(data_in[249]&H_in[3577])^(data_in[250]&H_in[3578])^(data_in[251]&H_in[3579])^(data_in[252]&H_in[3580])^(data_in[253]&H_in[3581])^(data_in[254]&H_in[3582])^(data_in[255]&H_in[3583]);
         data_out[14]<=data_out[14]^(data_in[0]&H_in[3584])^(data_in[1]&H_in[3585])^(data_in[2]&H_in[3586])^(data_in[3]&H_in[3587])^(data_in[4]&H_in[3588])^(data_in[5]&H_in[3589])^(data_in[6]&H_in[3590])^(data_in[7]&H_in[3591])^(data_in[8]&H_in[3592])^(data_in[9]&H_in[3593])^(data_in[10]&H_in[3594])^(data_in[11]&H_in[3595])^(data_in[12]&H_in[3596])^(data_in[13]&H_in[3597])^(data_in[14]&H_in[3598])^(data_in[15]&H_in[3599])^(data_in[16]&H_in[3600])^(data_in[17]&H_in[3601])^(data_in[18]&H_in[3602])^(data_in[19]&H_in[3603])^(data_in[20]&H_in[3604])^(data_in[21]&H_in[3605])^(data_in[22]&H_in[3606])^(data_in[23]&H_in[3607])^(data_in[24]&H_in[3608])^(data_in[25]&H_in[3609])^(data_in[26]&H_in[3610])^(data_in[27]&H_in[3611])^(data_in[28]&H_in[3612])^(data_in[29]&H_in[3613])^(data_in[30]&H_in[3614])^(data_in[31]&H_in[3615])^(data_in[32]&H_in[3616])^(data_in[33]&H_in[3617])^(data_in[34]&H_in[3618])^(data_in[35]&H_in[3619])^(data_in[36]&H_in[3620])^(data_in[37]&H_in[3621])^(data_in[38]&H_in[3622])^(data_in[39]&H_in[3623])^(data_in[40]&H_in[3624])^(data_in[41]&H_in[3625])^(data_in[42]&H_in[3626])^(data_in[43]&H_in[3627])^(data_in[44]&H_in[3628])^(data_in[45]&H_in[3629])^(data_in[46]&H_in[3630])^(data_in[47]&H_in[3631])^(data_in[48]&H_in[3632])^(data_in[49]&H_in[3633])^(data_in[50]&H_in[3634])^(data_in[51]&H_in[3635])^(data_in[52]&H_in[3636])^(data_in[53]&H_in[3637])^(data_in[54]&H_in[3638])^(data_in[55]&H_in[3639])^(data_in[56]&H_in[3640])^(data_in[57]&H_in[3641])^(data_in[58]&H_in[3642])^(data_in[59]&H_in[3643])^(data_in[60]&H_in[3644])^(data_in[61]&H_in[3645])^(data_in[62]&H_in[3646])^(data_in[63]&H_in[3647])^(data_in[64]&H_in[3648])^(data_in[65]&H_in[3649])^(data_in[66]&H_in[3650])^(data_in[67]&H_in[3651])^(data_in[68]&H_in[3652])^(data_in[69]&H_in[3653])^(data_in[70]&H_in[3654])^(data_in[71]&H_in[3655])^(data_in[72]&H_in[3656])^(data_in[73]&H_in[3657])^(data_in[74]&H_in[3658])^(data_in[75]&H_in[3659])^(data_in[76]&H_in[3660])^(data_in[77]&H_in[3661])^(data_in[78]&H_in[3662])^(data_in[79]&H_in[3663])^(data_in[80]&H_in[3664])^(data_in[81]&H_in[3665])^(data_in[82]&H_in[3666])^(data_in[83]&H_in[3667])^(data_in[84]&H_in[3668])^(data_in[85]&H_in[3669])^(data_in[86]&H_in[3670])^(data_in[87]&H_in[3671])^(data_in[88]&H_in[3672])^(data_in[89]&H_in[3673])^(data_in[90]&H_in[3674])^(data_in[91]&H_in[3675])^(data_in[92]&H_in[3676])^(data_in[93]&H_in[3677])^(data_in[94]&H_in[3678])^(data_in[95]&H_in[3679])^(data_in[96]&H_in[3680])^(data_in[97]&H_in[3681])^(data_in[98]&H_in[3682])^(data_in[99]&H_in[3683])^(data_in[100]&H_in[3684])^(data_in[101]&H_in[3685])^(data_in[102]&H_in[3686])^(data_in[103]&H_in[3687])^(data_in[104]&H_in[3688])^(data_in[105]&H_in[3689])^(data_in[106]&H_in[3690])^(data_in[107]&H_in[3691])^(data_in[108]&H_in[3692])^(data_in[109]&H_in[3693])^(data_in[110]&H_in[3694])^(data_in[111]&H_in[3695])^(data_in[112]&H_in[3696])^(data_in[113]&H_in[3697])^(data_in[114]&H_in[3698])^(data_in[115]&H_in[3699])^(data_in[116]&H_in[3700])^(data_in[117]&H_in[3701])^(data_in[118]&H_in[3702])^(data_in[119]&H_in[3703])^(data_in[120]&H_in[3704])^(data_in[121]&H_in[3705])^(data_in[122]&H_in[3706])^(data_in[123]&H_in[3707])^(data_in[124]&H_in[3708])^(data_in[125]&H_in[3709])^(data_in[126]&H_in[3710])^(data_in[127]&H_in[3711])^(data_in[128]&H_in[3712])^(data_in[129]&H_in[3713])^(data_in[130]&H_in[3714])^(data_in[131]&H_in[3715])^(data_in[132]&H_in[3716])^(data_in[133]&H_in[3717])^(data_in[134]&H_in[3718])^(data_in[135]&H_in[3719])^(data_in[136]&H_in[3720])^(data_in[137]&H_in[3721])^(data_in[138]&H_in[3722])^(data_in[139]&H_in[3723])^(data_in[140]&H_in[3724])^(data_in[141]&H_in[3725])^(data_in[142]&H_in[3726])^(data_in[143]&H_in[3727])^(data_in[144]&H_in[3728])^(data_in[145]&H_in[3729])^(data_in[146]&H_in[3730])^(data_in[147]&H_in[3731])^(data_in[148]&H_in[3732])^(data_in[149]&H_in[3733])^(data_in[150]&H_in[3734])^(data_in[151]&H_in[3735])^(data_in[152]&H_in[3736])^(data_in[153]&H_in[3737])^(data_in[154]&H_in[3738])^(data_in[155]&H_in[3739])^(data_in[156]&H_in[3740])^(data_in[157]&H_in[3741])^(data_in[158]&H_in[3742])^(data_in[159]&H_in[3743])^(data_in[160]&H_in[3744])^(data_in[161]&H_in[3745])^(data_in[162]&H_in[3746])^(data_in[163]&H_in[3747])^(data_in[164]&H_in[3748])^(data_in[165]&H_in[3749])^(data_in[166]&H_in[3750])^(data_in[167]&H_in[3751])^(data_in[168]&H_in[3752])^(data_in[169]&H_in[3753])^(data_in[170]&H_in[3754])^(data_in[171]&H_in[3755])^(data_in[172]&H_in[3756])^(data_in[173]&H_in[3757])^(data_in[174]&H_in[3758])^(data_in[175]&H_in[3759])^(data_in[176]&H_in[3760])^(data_in[177]&H_in[3761])^(data_in[178]&H_in[3762])^(data_in[179]&H_in[3763])^(data_in[180]&H_in[3764])^(data_in[181]&H_in[3765])^(data_in[182]&H_in[3766])^(data_in[183]&H_in[3767])^(data_in[184]&H_in[3768])^(data_in[185]&H_in[3769])^(data_in[186]&H_in[3770])^(data_in[187]&H_in[3771])^(data_in[188]&H_in[3772])^(data_in[189]&H_in[3773])^(data_in[190]&H_in[3774])^(data_in[191]&H_in[3775])^(data_in[192]&H_in[3776])^(data_in[193]&H_in[3777])^(data_in[194]&H_in[3778])^(data_in[195]&H_in[3779])^(data_in[196]&H_in[3780])^(data_in[197]&H_in[3781])^(data_in[198]&H_in[3782])^(data_in[199]&H_in[3783])^(data_in[200]&H_in[3784])^(data_in[201]&H_in[3785])^(data_in[202]&H_in[3786])^(data_in[203]&H_in[3787])^(data_in[204]&H_in[3788])^(data_in[205]&H_in[3789])^(data_in[206]&H_in[3790])^(data_in[207]&H_in[3791])^(data_in[208]&H_in[3792])^(data_in[209]&H_in[3793])^(data_in[210]&H_in[3794])^(data_in[211]&H_in[3795])^(data_in[212]&H_in[3796])^(data_in[213]&H_in[3797])^(data_in[214]&H_in[3798])^(data_in[215]&H_in[3799])^(data_in[216]&H_in[3800])^(data_in[217]&H_in[3801])^(data_in[218]&H_in[3802])^(data_in[219]&H_in[3803])^(data_in[220]&H_in[3804])^(data_in[221]&H_in[3805])^(data_in[222]&H_in[3806])^(data_in[223]&H_in[3807])^(data_in[224]&H_in[3808])^(data_in[225]&H_in[3809])^(data_in[226]&H_in[3810])^(data_in[227]&H_in[3811])^(data_in[228]&H_in[3812])^(data_in[229]&H_in[3813])^(data_in[230]&H_in[3814])^(data_in[231]&H_in[3815])^(data_in[232]&H_in[3816])^(data_in[233]&H_in[3817])^(data_in[234]&H_in[3818])^(data_in[235]&H_in[3819])^(data_in[236]&H_in[3820])^(data_in[237]&H_in[3821])^(data_in[238]&H_in[3822])^(data_in[239]&H_in[3823])^(data_in[240]&H_in[3824])^(data_in[241]&H_in[3825])^(data_in[242]&H_in[3826])^(data_in[243]&H_in[3827])^(data_in[244]&H_in[3828])^(data_in[245]&H_in[3829])^(data_in[246]&H_in[3830])^(data_in[247]&H_in[3831])^(data_in[248]&H_in[3832])^(data_in[249]&H_in[3833])^(data_in[250]&H_in[3834])^(data_in[251]&H_in[3835])^(data_in[252]&H_in[3836])^(data_in[253]&H_in[3837])^(data_in[254]&H_in[3838])^(data_in[255]&H_in[3839]);
         data_out[15]<=data_out[15]^(data_in[0]&H_in[3840])^(data_in[1]&H_in[3841])^(data_in[2]&H_in[3842])^(data_in[3]&H_in[3843])^(data_in[4]&H_in[3844])^(data_in[5]&H_in[3845])^(data_in[6]&H_in[3846])^(data_in[7]&H_in[3847])^(data_in[8]&H_in[3848])^(data_in[9]&H_in[3849])^(data_in[10]&H_in[3850])^(data_in[11]&H_in[3851])^(data_in[12]&H_in[3852])^(data_in[13]&H_in[3853])^(data_in[14]&H_in[3854])^(data_in[15]&H_in[3855])^(data_in[16]&H_in[3856])^(data_in[17]&H_in[3857])^(data_in[18]&H_in[3858])^(data_in[19]&H_in[3859])^(data_in[20]&H_in[3860])^(data_in[21]&H_in[3861])^(data_in[22]&H_in[3862])^(data_in[23]&H_in[3863])^(data_in[24]&H_in[3864])^(data_in[25]&H_in[3865])^(data_in[26]&H_in[3866])^(data_in[27]&H_in[3867])^(data_in[28]&H_in[3868])^(data_in[29]&H_in[3869])^(data_in[30]&H_in[3870])^(data_in[31]&H_in[3871])^(data_in[32]&H_in[3872])^(data_in[33]&H_in[3873])^(data_in[34]&H_in[3874])^(data_in[35]&H_in[3875])^(data_in[36]&H_in[3876])^(data_in[37]&H_in[3877])^(data_in[38]&H_in[3878])^(data_in[39]&H_in[3879])^(data_in[40]&H_in[3880])^(data_in[41]&H_in[3881])^(data_in[42]&H_in[3882])^(data_in[43]&H_in[3883])^(data_in[44]&H_in[3884])^(data_in[45]&H_in[3885])^(data_in[46]&H_in[3886])^(data_in[47]&H_in[3887])^(data_in[48]&H_in[3888])^(data_in[49]&H_in[3889])^(data_in[50]&H_in[3890])^(data_in[51]&H_in[3891])^(data_in[52]&H_in[3892])^(data_in[53]&H_in[3893])^(data_in[54]&H_in[3894])^(data_in[55]&H_in[3895])^(data_in[56]&H_in[3896])^(data_in[57]&H_in[3897])^(data_in[58]&H_in[3898])^(data_in[59]&H_in[3899])^(data_in[60]&H_in[3900])^(data_in[61]&H_in[3901])^(data_in[62]&H_in[3902])^(data_in[63]&H_in[3903])^(data_in[64]&H_in[3904])^(data_in[65]&H_in[3905])^(data_in[66]&H_in[3906])^(data_in[67]&H_in[3907])^(data_in[68]&H_in[3908])^(data_in[69]&H_in[3909])^(data_in[70]&H_in[3910])^(data_in[71]&H_in[3911])^(data_in[72]&H_in[3912])^(data_in[73]&H_in[3913])^(data_in[74]&H_in[3914])^(data_in[75]&H_in[3915])^(data_in[76]&H_in[3916])^(data_in[77]&H_in[3917])^(data_in[78]&H_in[3918])^(data_in[79]&H_in[3919])^(data_in[80]&H_in[3920])^(data_in[81]&H_in[3921])^(data_in[82]&H_in[3922])^(data_in[83]&H_in[3923])^(data_in[84]&H_in[3924])^(data_in[85]&H_in[3925])^(data_in[86]&H_in[3926])^(data_in[87]&H_in[3927])^(data_in[88]&H_in[3928])^(data_in[89]&H_in[3929])^(data_in[90]&H_in[3930])^(data_in[91]&H_in[3931])^(data_in[92]&H_in[3932])^(data_in[93]&H_in[3933])^(data_in[94]&H_in[3934])^(data_in[95]&H_in[3935])^(data_in[96]&H_in[3936])^(data_in[97]&H_in[3937])^(data_in[98]&H_in[3938])^(data_in[99]&H_in[3939])^(data_in[100]&H_in[3940])^(data_in[101]&H_in[3941])^(data_in[102]&H_in[3942])^(data_in[103]&H_in[3943])^(data_in[104]&H_in[3944])^(data_in[105]&H_in[3945])^(data_in[106]&H_in[3946])^(data_in[107]&H_in[3947])^(data_in[108]&H_in[3948])^(data_in[109]&H_in[3949])^(data_in[110]&H_in[3950])^(data_in[111]&H_in[3951])^(data_in[112]&H_in[3952])^(data_in[113]&H_in[3953])^(data_in[114]&H_in[3954])^(data_in[115]&H_in[3955])^(data_in[116]&H_in[3956])^(data_in[117]&H_in[3957])^(data_in[118]&H_in[3958])^(data_in[119]&H_in[3959])^(data_in[120]&H_in[3960])^(data_in[121]&H_in[3961])^(data_in[122]&H_in[3962])^(data_in[123]&H_in[3963])^(data_in[124]&H_in[3964])^(data_in[125]&H_in[3965])^(data_in[126]&H_in[3966])^(data_in[127]&H_in[3967])^(data_in[128]&H_in[3968])^(data_in[129]&H_in[3969])^(data_in[130]&H_in[3970])^(data_in[131]&H_in[3971])^(data_in[132]&H_in[3972])^(data_in[133]&H_in[3973])^(data_in[134]&H_in[3974])^(data_in[135]&H_in[3975])^(data_in[136]&H_in[3976])^(data_in[137]&H_in[3977])^(data_in[138]&H_in[3978])^(data_in[139]&H_in[3979])^(data_in[140]&H_in[3980])^(data_in[141]&H_in[3981])^(data_in[142]&H_in[3982])^(data_in[143]&H_in[3983])^(data_in[144]&H_in[3984])^(data_in[145]&H_in[3985])^(data_in[146]&H_in[3986])^(data_in[147]&H_in[3987])^(data_in[148]&H_in[3988])^(data_in[149]&H_in[3989])^(data_in[150]&H_in[3990])^(data_in[151]&H_in[3991])^(data_in[152]&H_in[3992])^(data_in[153]&H_in[3993])^(data_in[154]&H_in[3994])^(data_in[155]&H_in[3995])^(data_in[156]&H_in[3996])^(data_in[157]&H_in[3997])^(data_in[158]&H_in[3998])^(data_in[159]&H_in[3999])^(data_in[160]&H_in[4000])^(data_in[161]&H_in[4001])^(data_in[162]&H_in[4002])^(data_in[163]&H_in[4003])^(data_in[164]&H_in[4004])^(data_in[165]&H_in[4005])^(data_in[166]&H_in[4006])^(data_in[167]&H_in[4007])^(data_in[168]&H_in[4008])^(data_in[169]&H_in[4009])^(data_in[170]&H_in[4010])^(data_in[171]&H_in[4011])^(data_in[172]&H_in[4012])^(data_in[173]&H_in[4013])^(data_in[174]&H_in[4014])^(data_in[175]&H_in[4015])^(data_in[176]&H_in[4016])^(data_in[177]&H_in[4017])^(data_in[178]&H_in[4018])^(data_in[179]&H_in[4019])^(data_in[180]&H_in[4020])^(data_in[181]&H_in[4021])^(data_in[182]&H_in[4022])^(data_in[183]&H_in[4023])^(data_in[184]&H_in[4024])^(data_in[185]&H_in[4025])^(data_in[186]&H_in[4026])^(data_in[187]&H_in[4027])^(data_in[188]&H_in[4028])^(data_in[189]&H_in[4029])^(data_in[190]&H_in[4030])^(data_in[191]&H_in[4031])^(data_in[192]&H_in[4032])^(data_in[193]&H_in[4033])^(data_in[194]&H_in[4034])^(data_in[195]&H_in[4035])^(data_in[196]&H_in[4036])^(data_in[197]&H_in[4037])^(data_in[198]&H_in[4038])^(data_in[199]&H_in[4039])^(data_in[200]&H_in[4040])^(data_in[201]&H_in[4041])^(data_in[202]&H_in[4042])^(data_in[203]&H_in[4043])^(data_in[204]&H_in[4044])^(data_in[205]&H_in[4045])^(data_in[206]&H_in[4046])^(data_in[207]&H_in[4047])^(data_in[208]&H_in[4048])^(data_in[209]&H_in[4049])^(data_in[210]&H_in[4050])^(data_in[211]&H_in[4051])^(data_in[212]&H_in[4052])^(data_in[213]&H_in[4053])^(data_in[214]&H_in[4054])^(data_in[215]&H_in[4055])^(data_in[216]&H_in[4056])^(data_in[217]&H_in[4057])^(data_in[218]&H_in[4058])^(data_in[219]&H_in[4059])^(data_in[220]&H_in[4060])^(data_in[221]&H_in[4061])^(data_in[222]&H_in[4062])^(data_in[223]&H_in[4063])^(data_in[224]&H_in[4064])^(data_in[225]&H_in[4065])^(data_in[226]&H_in[4066])^(data_in[227]&H_in[4067])^(data_in[228]&H_in[4068])^(data_in[229]&H_in[4069])^(data_in[230]&H_in[4070])^(data_in[231]&H_in[4071])^(data_in[232]&H_in[4072])^(data_in[233]&H_in[4073])^(data_in[234]&H_in[4074])^(data_in[235]&H_in[4075])^(data_in[236]&H_in[4076])^(data_in[237]&H_in[4077])^(data_in[238]&H_in[4078])^(data_in[239]&H_in[4079])^(data_in[240]&H_in[4080])^(data_in[241]&H_in[4081])^(data_in[242]&H_in[4082])^(data_in[243]&H_in[4083])^(data_in[244]&H_in[4084])^(data_in[245]&H_in[4085])^(data_in[246]&H_in[4086])^(data_in[247]&H_in[4087])^(data_in[248]&H_in[4088])^(data_in[249]&H_in[4089])^(data_in[250]&H_in[4090])^(data_in[251]&H_in[4091])^(data_in[252]&H_in[4092])^(data_in[253]&H_in[4093])^(data_in[254]&H_in[4094])^(data_in[255]&H_in[4095]);

         end
         else begin 
             data_out <=data_out ;
         end
     end


    endmodule


